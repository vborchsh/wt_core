
`ifndef __WT_HEADER__
`define __WT_HEADER__

//--------------------------------------------------------------------------------------------------------
// File connection
//--------------------------------------------------------------------------------------------------------

//
`include "./../rtl/wt_common/wt_fir.sv"
`include "./../rtl/idwt_core.sv"
`include "./../rtl/dwt_core.sv"

//--------------------------------------------------------------------------------------------------------
// Parameters
//--------------------------------------------------------------------------------------------------------


`endif

