
module tb_wt_fir;
  // ******************************************
  // CLOCK GENERATOR***************************
  timeunit 1ns;
  timeprecision 1ns;

  bit  clk;
  initial begin
    forever #1 clk = ~clk;
  end
  // ******************************************
  // ******************************************
  
  //--------------------------------------------------------------------------------------------------
  // Declaration parameters
  //--------------------------------------------------------------------------------------------------

  localparam int pWIDTH = 12;
  localparam int pORDER = 12;
  localparam int cCOEFS [pORDER] = '{-5,  19,  2,  -130,  112,  399,  -532,  -927,  1291,  3076,  2025,  456};
 
  //--------------------------------------------------------------------------------------------------
  // Declaration variables
  //--------------------------------------------------------------------------------------------------
  
  logic           [7:0] arr          [128];
  logic           [3:0] cnt_ena      ;
  logic                 clk_ena      ;
  //
  logic                 fir__iclk    ;
  logic                 fir__iclk_ena;
  logic                 fir__irst    ;
  logic                 fir__iena    ;
  logic    [pWIDTH-1:0] fir__idat    ;
  logic                 fir__oena    ;
  logic  [2*pWIDTH-1:0] fir__odat    ;

  //--------------------------------------------------------------------------------------------------
  // Initialization
  //--------------------------------------------------------------------------------------------------

  initial begin
    for (int i = 0; i < $size(arr); i++) begin
      arr[i] = 0;
      //arr[i] = $urandom_range(0, 64);
      //arr[i] = i;
    end
    //
    arr[64] = '1;
  end
  
  //--------------------------------------------------------------------------------------------------
  // BODY
  //--------------------------------------------------------------------------------------------------

  always@(posedge clk) begin
    cnt_ena <= cnt_ena + 1'b1;
    clk_ena <= &cnt_ena;
  end
  // Main thread
  initial begin
    
  end

  //--------------------------------------------------------------------------------------------------
  // Modules
  //--------------------------------------------------------------------------------------------------

  wt_fir
  #(
    . pWIDTH     (pWIDTH        ) ,
    . pORDER     (pORDER        ) ,
    . cCOEFS     (cCOEFS        )
  )
  fir__
  (
    . iclk       (clk           ) ,
    . iclk_ena   (clk_ena       ) ,
    . irst       (fir__irst     ) ,
    . iena       (fir__iena     ) ,
    . idat       (fir__idat     ) ,
    . oena       (fir__oena     ) ,
    . odat       (fir__odat     )
  );

endmodule
