
`ifndef __WT_HEADER__
`define __WT_HEADER__

//--------------------------------------------------------------------------------------------------------
// File connection
//--------------------------------------------------------------------------------------------------------

//
`include "./../rtl/wt_common/wt_fir.sv"

//--------------------------------------------------------------------------------------------------------
// Parameters
//--------------------------------------------------------------------------------------------------------


`endif

