
`ifndef __WT_WAVELETS__
`define __WT_WAVELETS__

localparam real pHAAR_Lo_D [2] = '{0.707106781186547570000000,0.707106781186547570000000};
localparam real pHAAR_Lo_R [2] = '{0.707106781186547570000000,0.707106781186547570000000};
localparam real pHAAR_Hi_D [2] = '{-0.707106781186547570000000,0.707106781186547570000000};
localparam real pHAAR_Hi_R [2] = '{0.707106781186547570000000,-0.707106781186547570000000};

localparam real pDB1_Lo_D [2] = '{0.707106781186547570000000,0.707106781186547570000000};
localparam real pDB1_Lo_R [2] = '{0.707106781186547570000000,0.707106781186547570000000};
localparam real pDB1_Hi_D [2] = '{-0.707106781186547570000000,0.707106781186547570000000};
localparam real pDB1_Hi_R [2] = '{0.707106781186547570000000,-0.707106781186547570000000};

localparam real pDB2_Lo_D [4] = '{-0.129409522550921450000000,0.224143868041857350000000,0.836516303737468990000000,0.482962913144690250000000};
localparam real pDB2_Lo_R [4] = '{0.482962913144690250000000,0.836516303737468990000000,0.224143868041857350000000,-0.129409522550921450000000};
localparam real pDB2_Hi_D [4] = '{-0.482962913144690250000000,0.836516303737468990000000,-0.224143868041857350000000,-0.129409522550921450000000};
localparam real pDB2_Hi_R [4] = '{-0.129409522550921450000000,-0.224143868041857350000000,0.836516303737468990000000,-0.482962913144690250000000};

localparam real pDB3_Lo_D [6] = '{0.035226291882100656000000,-0.085441273882241486000000,-0.135011020010390840000000,0.459877502119331320000000,0.806891509313338750000000,0.332670552950956880000000};
localparam real pDB3_Lo_R [6] = '{0.332670552950956880000000,0.806891509313338750000000,0.459877502119331320000000,-0.135011020010390840000000,-0.085441273882241486000000,0.035226291882100656000000};
localparam real pDB3_Hi_D [6] = '{-0.332670552950956880000000,0.806891509313338750000000,-0.459877502119331320000000,-0.135011020010390840000000,0.085441273882241486000000,0.035226291882100656000000};
localparam real pDB3_Hi_R [6] = '{0.035226291882100656000000,0.085441273882241486000000,-0.135011020010390840000000,-0.459877502119331320000000,0.806891509313338750000000,-0.332670552950956880000000};

localparam real pDB4_Lo_D [8] = '{-0.010597401784997278000000,0.032883011666982945000000,0.030841381835986965000000,-0.187034811718881140000000,-0.027983769416983849000000,0.630880767929590360000000,0.714846570552541530000000,0.230377813308855230000000};
localparam real pDB4_Lo_R [8] = '{0.230377813308855230000000,0.714846570552541530000000,0.630880767929590360000000,-0.027983769416983849000000,-0.187034811718881140000000,0.030841381835986965000000,0.032883011666982945000000,-0.010597401784997278000000};
localparam real pDB4_Hi_D [8] = '{-0.230377813308855230000000,0.714846570552541530000000,-0.630880767929590360000000,-0.027983769416983849000000,0.187034811718881140000000,0.030841381835986965000000,-0.032883011666982945000000,-0.010597401784997278000000};
localparam real pDB4_Hi_R [8] = '{-0.010597401784997278000000,-0.032883011666982945000000,0.030841381835986965000000,0.187034811718881140000000,-0.027983769416983849000000,-0.630880767929590360000000,0.714846570552541530000000,-0.230377813308855230000000};

localparam real pDB5_Lo_D [10] = '{0.003335725285001549200000,-0.012580751999015526000000,-0.006241490213011705200000,0.077571493840065148000000,-0.032244869585029520000000,-0.242294887066190150000000,0.138428145901103420000000,0.724308528438574410000000,0.603829269797472870000000,0.160102397974125010000000};
localparam real pDB5_Lo_R [10] = '{0.160102397974125010000000,0.603829269797472870000000,0.724308528438574410000000,0.138428145901103420000000,-0.242294887066190150000000,-0.032244869585029520000000,0.077571493840065148000000,-0.006241490213011705200000,-0.012580751999015526000000,0.003335725285001549200000};
localparam real pDB5_Hi_D [10] = '{-0.160102397974125010000000,0.603829269797472870000000,-0.724308528438574410000000,0.138428145901103420000000,0.242294887066190150000000,-0.032244869585029520000000,-0.077571493840065148000000,-0.006241490213011705200000,0.012580751999015526000000,0.003335725285001549200000};
localparam real pDB5_Hi_R [10] = '{0.003335725285001549200000,0.012580751999015526000000,-0.006241490213011705200000,-0.077571493840065148000000,-0.032244869585029520000000,0.242294887066190150000000,0.138428145901103420000000,-0.724308528438574410000000,0.603829269797472870000000,-0.160102397974125010000000};

localparam real pDB6_Lo_D [12] = '{-0.001077301084995579900000,0.004777257511010651400000,0.000553842200993801600000,-0.031582039318031156000000,0.027522865530016288000000,0.097501605587079362000000,-0.129766867567095630000000,-0.226264693965169130000000,0.315250351709243200000000,0.751133908021577530000000,0.494623890398385390000000,0.111540743350080170000000};
localparam real pDB6_Lo_R [12] = '{0.111540743350080170000000,0.494623890398385390000000,0.751133908021577530000000,0.315250351709243200000000,-0.226264693965169130000000,-0.129766867567095630000000,0.097501605587079362000000,0.027522865530016288000000,-0.031582039318031156000000,0.000553842200993801600000,0.004777257511010651400000,-0.001077301084995579900000};
localparam real pDB6_Hi_D [12] = '{-0.111540743350080170000000,0.494623890398385390000000,-0.751133908021577530000000,0.315250351709243200000000,0.226264693965169130000000,-0.129766867567095630000000,-0.097501605587079362000000,0.027522865530016288000000,0.031582039318031156000000,0.000553842200993801600000,-0.004777257511010651400000,-0.001077301084995579900000};
localparam real pDB6_Hi_R [12] = '{-0.001077301084995579900000,-0.004777257511010651400000,0.000553842200993801600000,0.031582039318031156000000,0.027522865530016288000000,-0.097501605587079362000000,-0.129766867567095630000000,0.226264693965169130000000,0.315250351709243200000000,-0.751133908021577530000000,0.494623890398385390000000,-0.111540743350080170000000};

localparam real pDB7_Lo_D [14] = '{0.000353713800001039880000,-0.001801640703999832800000,0.000429577973004702740000,0.012550998556013784000000,-0.016574541631015620000000,-0.038029936935034633000000,0.080612609151065898000000,0.071309219267050042000000,-0.224036184994165720000000,-0.143906003929106270000000,0.469782287405358600000000,0.729132090846555060000000,0.396539319482305750000000,0.077852054085062364000000};
localparam real pDB7_Lo_R [14] = '{0.077852054085062364000000,0.396539319482305750000000,0.729132090846555060000000,0.469782287405358600000000,-0.143906003929106270000000,-0.224036184994165720000000,0.071309219267050042000000,0.080612609151065898000000,-0.038029936935034633000000,-0.016574541631015620000000,0.012550998556013784000000,0.000429577973004702740000,-0.001801640703999832800000,0.000353713800001039880000};
localparam real pDB7_Hi_D [14] = '{-0.077852054085062364000000,0.396539319482305750000000,-0.729132090846555060000000,0.469782287405358600000000,0.143906003929106270000000,-0.224036184994165720000000,-0.071309219267050042000000,0.080612609151065898000000,0.038029936935034633000000,-0.016574541631015620000000,-0.012550998556013784000000,0.000429577973004702740000,0.001801640703999832800000,0.000353713800001039880000};
localparam real pDB7_Hi_R [14] = '{0.000353713800001039880000,0.001801640703999832800000,0.000429577973004702740000,-0.012550998556013784000000,-0.016574541631015620000000,0.038029936935034633000000,0.080612609151065898000000,-0.071309219267050042000000,-0.224036184994165720000000,0.143906003929106270000000,0.469782287405358600000000,-0.729132090846555060000000,0.396539319482305750000000,-0.077852054085062364000000};

localparam real pDB8_Lo_D [16] = '{-0.000117476784002281920000,0.000675449405998556770000,-0.000391740372995977110000,-0.004870352993010660300000,0.008746094047015654700000,0.013981027917015516000000,-0.044088253931064719000000,-0.017369301002022108000000,0.128747426620186010000000,0.000472484573997972540000,-0.284015542962428090000000,-0.015829105256023893000000,0.585354683654869090000000,0.675630736298012850000000,0.312871590914465920000000,0.054415842243081609000000};
localparam real pDB8_Lo_R [16] = '{0.054415842243081609000000,0.312871590914465920000000,0.675630736298012850000000,0.585354683654869090000000,-0.015829105256023893000000,-0.284015542962428090000000,0.000472484573997972540000,0.128747426620186010000000,-0.017369301002022108000000,-0.044088253931064719000000,0.013981027917015516000000,0.008746094047015654700000,-0.004870352993010660300000,-0.000391740372995977110000,0.000675449405998556770000,-0.000117476784002281920000};
localparam real pDB8_Hi_D [16] = '{-0.054415842243081609000000,0.312871590914465920000000,-0.675630736298012850000000,0.585354683654869090000000,0.015829105256023893000000,-0.284015542962428090000000,-0.000472484573997972540000,0.128747426620186010000000,0.017369301002022108000000,-0.044088253931064719000000,-0.013981027917015516000000,0.008746094047015654700000,0.004870352993010660300000,-0.000391740372995977110000,-0.000675449405998556770000,-0.000117476784002281920000};
localparam real pDB8_Hi_R [16] = '{-0.000117476784002281920000,-0.000675449405998556770000,-0.000391740372995977110000,0.004870352993010660300000,0.008746094047015654700000,-0.013981027917015516000000,-0.044088253931064719000000,0.017369301002022108000000,0.128747426620186010000000,-0.000472484573997972540000,-0.284015542962428090000000,0.015829105256023893000000,0.585354683654869090000000,-0.675630736298012850000000,0.312871590914465920000000,-0.054415842243081609000000};

localparam real pDB9_Lo_D [18] = '{0.000039347319995026124000,-0.000251963188998178880000,0.000230385763995412880000,0.001847646882961126800000,-0.004281503681904722700000,-0.004723204757894831000000,0.022361662123515244000000,0.000250947114991938450000,-0.067632829059523988000000,0.030725681478322865000000,0.148540749334760080000000,-0.096840783220879037000000,-0.293273783272586850000000,0.133197385822088950000000,0.657288078036638910000000,0.604823123676778600000000,0.243834674637667280000000,0.038077947363167282000000};
localparam real pDB9_Lo_R [18] = '{0.038077947363167282000000,0.243834674637667280000000,0.604823123676778600000000,0.657288078036638910000000,0.133197385822088950000000,-0.293273783272586850000000,-0.096840783220879037000000,0.148540749334760080000000,0.030725681478322865000000,-0.067632829059523988000000,0.000250947114991938450000,0.022361662123515244000000,-0.004723204757894831000000,-0.004281503681904722700000,0.001847646882961126800000,0.000230385763995412880000,-0.000251963188998178880000,0.000039347319995026124000};
localparam real pDB9_Hi_D [18] = '{-0.038077947363167282000000,0.243834674637667280000000,-0.604823123676778600000000,0.657288078036638910000000,-0.133197385822088950000000,-0.293273783272586850000000,0.096840783220879037000000,0.148540749334760080000000,-0.030725681478322865000000,-0.067632829059523988000000,-0.000250947114991938450000,0.022361662123515244000000,0.004723204757894831000000,-0.004281503681904722700000,-0.001847646882961126800000,0.000230385763995412880000,0.000251963188998178880000,0.000039347319995026124000};
localparam real pDB9_Hi_R [18] = '{0.000039347319995026124000,0.000251963188998178880000,0.000230385763995412880000,-0.001847646882961126800000,-0.004281503681904722700000,0.004723204757894831000000,0.022361662123515244000000,-0.000250947114991938450000,-0.067632829059523988000000,-0.030725681478322865000000,0.148540749334760080000000,0.096840783220879037000000,-0.293273783272586850000000,-0.133197385822088950000000,0.657288078036638910000000,-0.604823123676778600000000,0.243834674637667280000000,-0.038077947363167282000000};

localparam real pDB10_Lo_D [20] = '{-0.000013264203002354869000,0.000093588670001089845000,-0.000116466854994386200000,-0.000685856695004682480000,0.001992405294990849900000,0.001395351746994079800000,-0.010733175482979604000000,0.003606553566988394400000,0.033212674058933238000000,-0.029457536821945671000000,-0.071394147165860775000000,0.093057364603806592000000,0.127369340335742650000000,-0.195946274376596650000000,-0.249846424326488650000000,0.281172343660426480000000,0.688459039452592130000000,0.527201188930919830000000,0.188176800077621330000000,0.026670057900950818000000};
localparam real pDB10_Lo_R [20] = '{0.026670057900950818000000,0.188176800077621330000000,0.527201188930919830000000,0.688459039452592130000000,0.281172343660426480000000,-0.249846424326488650000000,-0.195946274376596650000000,0.127369340335742650000000,0.093057364603806592000000,-0.071394147165860775000000,-0.029457536821945671000000,0.033212674058933238000000,0.003606553566988394400000,-0.010733175482979604000000,0.001395351746994079800000,0.001992405294990849900000,-0.000685856695004682480000,-0.000116466854994386200000,0.000093588670001089845000,-0.000013264203002354869000};
localparam real pDB10_Hi_D [20] = '{-0.026670057900950818000000,0.188176800077621330000000,-0.527201188930919830000000,0.688459039452592130000000,-0.281172343660426480000000,-0.249846424326488650000000,0.195946274376596650000000,0.127369340335742650000000,-0.093057364603806592000000,-0.071394147165860775000000,0.029457536821945671000000,0.033212674058933238000000,-0.003606553566988394400000,-0.010733175482979604000000,-0.001395351746994079800000,0.001992405294990849900000,0.000685856695004682480000,-0.000116466854994386200000,-0.000093588670001089845000,-0.000013264203002354869000};
localparam real pDB10_Hi_R [20] = '{-0.000013264203002354869000,-0.000093588670001089845000,-0.000116466854994386200000,0.000685856695004682480000,0.001992405294990849900000,-0.001395351746994079800000,-0.010733175482979604000000,-0.003606553566988394400000,0.033212674058933238000000,0.029457536821945671000000,-0.071394147165860775000000,-0.093057364603806592000000,0.127369340335742650000000,0.195946274376596650000000,-0.249846424326488650000000,-0.281172343660426480000000,0.688459039452592130000000,-0.527201188930919830000000,0.188176800077621330000000,-0.026670057900950818000000};

localparam real pDB11_Lo_D [22] = '{0.000004494274277236586500,-0.000034634984186985538000,0.000054439074699369044000,0.000249152523552826240000,-0.000893023250666285530000,-0.000308592858815184390000,0.004928417656059012700000,-0.003340858873014710400000,-0.015364820906202272000000,0.020840904360180473000000,0.031335090219044910000000,-0.066438785695028771000000,-0.046479955116688516000000,0.149812012466376380000000,0.066043588196680117000000,-0.274230846817953680000000,-0.162275245027493710000000,0.411964368947913720000000,0.685686774916211110000000,0.449899764356052110000000,0.144067021150626700000000,0.018694297761471367000000};
localparam real pDB11_Lo_R [22] = '{0.018694297761471367000000,0.144067021150626700000000,0.449899764356052110000000,0.685686774916211110000000,0.411964368947913720000000,-0.162275245027493710000000,-0.274230846817953680000000,0.066043588196680117000000,0.149812012466376380000000,-0.046479955116688516000000,-0.066438785695028771000000,0.031335090219044910000000,0.020840904360180473000000,-0.015364820906202272000000,-0.003340858873014710400000,0.004928417656059012700000,-0.000308592858815184390000,-0.000893023250666285530000,0.000249152523552826240000,0.000054439074699369044000,-0.000034634984186985538000,0.000004494274277236586500};
localparam real pDB11_Hi_D [22] = '{-0.018694297761471367000000,0.144067021150626700000000,-0.449899764356052110000000,0.685686774916211110000000,-0.411964368947913720000000,-0.162275245027493710000000,0.274230846817953680000000,0.066043588196680117000000,-0.149812012466376380000000,-0.046479955116688516000000,0.066438785695028771000000,0.031335090219044910000000,-0.020840904360180473000000,-0.015364820906202272000000,0.003340858873014710400000,0.004928417656059012700000,0.000308592858815184390000,-0.000893023250666285530000,-0.000249152523552826240000,0.000054439074699369044000,0.000034634984186985538000,0.000004494274277236586500};
localparam real pDB11_Hi_R [22] = '{0.000004494274277236586500,0.000034634984186985538000,0.000054439074699369044000,-0.000249152523552826240000,-0.000893023250666285530000,0.000308592858815184390000,0.004928417656059012700000,0.003340858873014710400000,-0.015364820906202272000000,-0.020840904360180473000000,0.031335090219044910000000,0.066438785695028771000000,-0.046479955116688516000000,-0.149812012466376380000000,0.066043588196680117000000,0.274230846817953680000000,-0.162275245027493710000000,-0.411964368947913720000000,0.685686774916211110000000,-0.449899764356052110000000,0.144067021150626700000000,-0.018694297761471367000000};

localparam real pDB12_Lo_D [24] = '{-0.000001529071758068568700,0.000012776952219380249000,-0.000024241545757031649000,-0.000088504109208206976000,0.000388653062820950410000,0.000006545128212521341700,-0.002179503618627852700000,0.002248607240995142800000,0.006711499008795106200000,-0.012840825198302545000000,-0.012218649069750715000000,0.041546277495083647000000,0.010849130255819399000000,-0.096432120096515805000000,0.005359569674345064800000,0.182478605927578170000000,-0.023779257256078486000000,-0.316178453752803850000000,-0.044763885653780866000000,0.515886478427832420000000,0.657198722579330650000000,0.377355135214226530000000,0.109566272821189220000000,0.013112257957230007000000};
localparam real pDB12_Lo_R [24] = '{0.013112257957230007000000,0.109566272821189220000000,0.377355135214226530000000,0.657198722579330650000000,0.515886478427832420000000,-0.044763885653780866000000,-0.316178453752803850000000,-0.023779257256078486000000,0.182478605927578170000000,0.005359569674345064800000,-0.096432120096515805000000,0.010849130255819399000000,0.041546277495083647000000,-0.012218649069750715000000,-0.012840825198302545000000,0.006711499008795106200000,0.002248607240995142800000,-0.002179503618627852700000,0.000006545128212521341700,0.000388653062820950410000,-0.000088504109208206976000,-0.000024241545757031649000,0.000012776952219380249000,-0.000001529071758068568700};
localparam real pDB12_Hi_D [24] = '{-0.013112257957230007000000,0.109566272821189220000000,-0.377355135214226530000000,0.657198722579330650000000,-0.515886478427832420000000,-0.044763885653780866000000,0.316178453752803850000000,-0.023779257256078486000000,-0.182478605927578170000000,0.005359569674345064800000,0.096432120096515805000000,0.010849130255819399000000,-0.041546277495083647000000,-0.012218649069750715000000,0.012840825198302545000000,0.006711499008795106200000,-0.002248607240995142800000,-0.002179503618627852700000,-0.000006545128212521341700,0.000388653062820950410000,0.000088504109208206976000,-0.000024241545757031649000,-0.000012776952219380249000,-0.000001529071758068568700};
localparam real pDB12_Hi_R [24] = '{-0.000001529071758068568700,-0.000012776952219380249000,-0.000024241545757031649000,0.000088504109208206976000,0.000388653062820950410000,-0.000006545128212521341700,-0.002179503618627852700000,-0.002248607240995142800000,0.006711499008795106200000,0.012840825198302545000000,-0.012218649069750715000000,-0.041546277495083647000000,0.010849130255819399000000,0.096432120096515805000000,0.005359569674345064800000,-0.182478605927578170000000,-0.023779257256078486000000,0.316178453752803850000000,-0.044763885653780866000000,-0.515886478427832420000000,0.657198722579330650000000,-0.377355135214226530000000,0.109566272821189220000000,-0.013112257957230007000000};

localparam real pDB13_Lo_D [26] = '{0.000000522003509845487390,-0.000004700416479360869200,0.000010441930571408100000,0.000030678537579325632000,-0.000165128988556502670000,0.000049251525126301336000,0.000932326130867286110000,-0.001315673911892272500000,-0.002761911234656847000000,0.007255589401617457000000,0.003923941448796887000000,-0.023831420710324711000000,0.002379972254058007900000,0.056139477100282859000000,-0.026488406475344117000000,-0.105807618187935020000000,0.072948933656776738000000,0.179476079429340050000000,-0.124576730750814990000000,-0.314972907711388360000000,0.086985726179647921000000,0.588889570431220140000000,0.611055851158788800000000,0.311996322160438600000000,0.082861243872902904000000,0.009202133538962382900000};
localparam real pDB13_Lo_R [26] = '{0.009202133538962382900000,0.082861243872902904000000,0.311996322160438600000000,0.611055851158788800000000,0.588889570431220140000000,0.086985726179647921000000,-0.314972907711388360000000,-0.124576730750814990000000,0.179476079429340050000000,0.072948933656776738000000,-0.105807618187935020000000,-0.026488406475344117000000,0.056139477100282859000000,0.002379972254058007900000,-0.023831420710324711000000,0.003923941448796887000000,0.007255589401617457000000,-0.002761911234656847000000,-0.001315673911892272500000,0.000932326130867286110000,0.000049251525126301336000,-0.000165128988556502670000,0.000030678537579325632000,0.000010441930571408100000,-0.000004700416479360869200,0.000000522003509845487390};
localparam real pDB13_Hi_D [26] = '{-0.009202133538962382900000,0.082861243872902904000000,-0.311996322160438600000000,0.611055851158788800000000,-0.588889570431220140000000,0.086985726179647921000000,0.314972907711388360000000,-0.124576730750814990000000,-0.179476079429340050000000,0.072948933656776738000000,0.105807618187935020000000,-0.026488406475344117000000,-0.056139477100282859000000,0.002379972254058007900000,0.023831420710324711000000,0.003923941448796887000000,-0.007255589401617457000000,-0.002761911234656847000000,0.001315673911892272500000,0.000932326130867286110000,-0.000049251525126301336000,-0.000165128988556502670000,-0.000030678537579325632000,0.000010441930571408100000,0.000004700416479360869200,0.000000522003509845487390};
localparam real pDB13_Hi_R [26] = '{0.000000522003509845487390,0.000004700416479360869200,0.000010441930571408100000,-0.000030678537579325632000,-0.000165128988556502670000,-0.000049251525126301336000,0.000932326130867286110000,0.001315673911892272500000,-0.002761911234656847000000,-0.007255589401617457000000,0.003923941448796887000000,0.023831420710324711000000,0.002379972254058007900000,-0.056139477100282859000000,-0.026488406475344117000000,0.105807618187935020000000,0.072948933656776738000000,-0.179476079429340050000000,-0.124576730750814990000000,0.314972907711388360000000,0.086985726179647921000000,-0.588889570431220140000000,0.611055851158788800000000,-0.311996322160438600000000,0.082861243872902904000000,-0.009202133538962382900000};

localparam real pDB14_Lo_D [28] = '{-0.000000178713996831074690,0.000001724994675367209800,-0.000004389704901779908500,-0.000010337209184567203000,0.000068755042526951268000,-0.000041777245770358305000,-0.000386831947312819410000,0.000708021154235258220000,0.001061691085606193200000,-0.003849638868021481800000,-0.000746218989269076040000,0.012789493266329202000000,-0.005615049530348897200000,-0.030185351540359097000000,0.026981408307948696000000,0.055237126259266384000000,-0.071548955503937847000000,-0.086748411568055253000000,0.139989016584486010000000,0.138395213864811380000000,-0.218033529993172850000000,-0.271688552278643360000000,0.218670687758836080000000,0.631187849104643320000000,0.554305617940705760000000,0.254850267792534890000000,0.062364758849377734000000,0.006461153460085754900000};
localparam real pDB14_Lo_R [28] = '{0.006461153460085754900000,0.062364758849377734000000,0.254850267792534890000000,0.554305617940705760000000,0.631187849104643320000000,0.218670687758836080000000,-0.271688552278643360000000,-0.218033529993172850000000,0.138395213864811380000000,0.139989016584486010000000,-0.086748411568055253000000,-0.071548955503937847000000,0.055237126259266384000000,0.026981408307948696000000,-0.030185351540359097000000,-0.005615049530348897200000,0.012789493266329202000000,-0.000746218989269076040000,-0.003849638868021481800000,0.001061691085606193200000,0.000708021154235258220000,-0.000386831947312819410000,-0.000041777245770358305000,0.000068755042526951268000,-0.000010337209184567203000,-0.000004389704901779908500,0.000001724994675367209800,-0.000000178713996831074690};
localparam real pDB14_Hi_D [28] = '{-0.006461153460085754900000,0.062364758849377734000000,-0.254850267792534890000000,0.554305617940705760000000,-0.631187849104643320000000,0.218670687758836080000000,0.271688552278643360000000,-0.218033529993172850000000,-0.138395213864811380000000,0.139989016584486010000000,0.086748411568055253000000,-0.071548955503937847000000,-0.055237126259266384000000,0.026981408307948696000000,0.030185351540359097000000,-0.005615049530348897200000,-0.012789493266329202000000,-0.000746218989269076040000,0.003849638868021481800000,0.001061691085606193200000,-0.000708021154235258220000,-0.000386831947312819410000,0.000041777245770358305000,0.000068755042526951268000,0.000010337209184567203000,-0.000004389704901779908500,-0.000001724994675367209800,-0.000000178713996831074690};
localparam real pDB14_Hi_R [28] = '{-0.000000178713996831074690,-0.000001724994675367209800,-0.000004389704901779908500,0.000010337209184567203000,0.000068755042526951268000,0.000041777245770358305000,-0.000386831947312819410000,-0.000708021154235258220000,0.001061691085606193200000,0.003849638868021481800000,-0.000746218989269076040000,-0.012789493266329202000000,-0.005615049530348897200000,0.030185351540359097000000,0.026981408307948696000000,-0.055237126259266384000000,-0.071548955503937847000000,0.086748411568055253000000,0.139989016584486010000000,-0.138395213864811380000000,-0.218033529993172850000000,0.271688552278643360000000,0.218670687758836080000000,-0.631187849104643320000000,0.554305617940705760000000,-0.254850267792534890000000,0.062364758849377734000000,-0.006461153460085754900000};

localparam real pDB15_Lo_D [30] = '{0.000000061333599133061239,-0.000000631688232588204250,0.000001811270407940691500,0.000003362987181737829000,-0.000028133296266049179000,0.000025792699155321555000,0.000155896489920613560000,-0.000359565244362451610000,-0.000373482354137428110000,0.001943323980382986200000,-0.000241756490760457130000,-0.006487734560315418400000,0.005101000360405317200000,0.015083918027827766000000,-0.020810050169709247000000,-0.025767007328454807000000,0.054780550584508134000000,0.033877143923517400000000,-0.111120936037230560000000,-0.039666176555795317000000,0.190146714007121350000000,0.065282952848758319000000,-0.288882596566999720000000,-0.193204139609167270000000,0.339002535454748570000000,0.645813140357463840000000,0.492631771708170410000000,0.206023863987008670000000,0.046743394892769220000000,0.004538537361579184600000};
localparam real pDB15_Lo_R [30] = '{0.004538537361579184600000,0.046743394892769220000000,0.206023863987008670000000,0.492631771708170410000000,0.645813140357463840000000,0.339002535454748570000000,-0.193204139609167270000000,-0.288882596566999720000000,0.065282952848758319000000,0.190146714007121350000000,-0.039666176555795317000000,-0.111120936037230560000000,0.033877143923517400000000,0.054780550584508134000000,-0.025767007328454807000000,-0.020810050169709247000000,0.015083918027827766000000,0.005101000360405317200000,-0.006487734560315418400000,-0.000241756490760457130000,0.001943323980382986200000,-0.000373482354137428110000,-0.000359565244362451610000,0.000155896489920613560000,0.000025792699155321555000,-0.000028133296266049179000,0.000003362987181737829000,0.000001811270407940691500,-0.000000631688232588204250,0.000000061333599133061239};
localparam real pDB15_Hi_D [30] = '{-0.004538537361579184600000,0.046743394892769220000000,-0.206023863987008670000000,0.492631771708170410000000,-0.645813140357463840000000,0.339002535454748570000000,0.193204139609167270000000,-0.288882596566999720000000,-0.065282952848758319000000,0.190146714007121350000000,0.039666176555795317000000,-0.111120936037230560000000,-0.033877143923517400000000,0.054780550584508134000000,0.025767007328454807000000,-0.020810050169709247000000,-0.015083918027827766000000,0.005101000360405317200000,0.006487734560315418400000,-0.000241756490760457130000,-0.001943323980382986200000,-0.000373482354137428110000,0.000359565244362451610000,0.000155896489920613560000,-0.000025792699155321555000,-0.000028133296266049179000,-0.000003362987181737829000,0.000001811270407940691500,0.000000631688232588204250,0.000000061333599133061239};
localparam real pDB15_Hi_R [30] = '{0.000000061333599133061239,0.000000631688232588204250,0.000001811270407940691500,-0.000003362987181737829000,-0.000028133296266049179000,-0.000025792699155321555000,0.000155896489920613560000,0.000359565244362451610000,-0.000373482354137428110000,-0.001943323980382986200000,-0.000241756490760457130000,0.006487734560315418400000,0.005101000360405317200000,-0.015083918027827766000000,-0.020810050169709247000000,0.025767007328454807000000,0.054780550584508134000000,-0.033877143923517400000000,-0.111120936037230560000000,0.039666176555795317000000,0.190146714007121350000000,-0.065282952848758319000000,-0.288882596566999720000000,0.193204139609167270000000,0.339002535454748570000000,-0.645813140357463840000000,0.492631771708170410000000,-0.206023863987008670000000,0.046743394892769220000000,-0.004538537361579184600000};

localparam real pDB16_Lo_D [32] = '{-0.000000021093396301004384,0.000000230878408685722150,-0.000000736365678545024900,-0.000001043571342311495000,0.000011336608661274467000,-0.000013945668988208811000,-0.000061035966214111162000,0.000174787245225280790000,0.000114241520038639420000,-0.000941021749359573200000,0.000407896980849087590000,0.003128023381203260100000,-0.003644279621506338400000,-0.006990014563432881200000,0.013993768859792647000000,0.010297659640913849000000,-0.036888397691750965000000,-0.007588974368841774000000,0.075924236044333640000000,-0.006239722752369098900000,-0.132388305563687660000000,0.027340263752781480000000,0.211190693947099300000000,-0.027918208133030944000000,-0.327063310527889450000000,-0.089751089402492351000000,0.440290256886286200000000,0.637356332083695460000000,0.430312722845942080000000,0.165064283488829620000000,0.034907714323668397000000,0.003189220925347287500000};
localparam real pDB16_Lo_R [32] = '{0.003189220925347287500000,0.034907714323668397000000,0.165064283488829620000000,0.430312722845942080000000,0.637356332083695460000000,0.440290256886286200000000,-0.089751089402492351000000,-0.327063310527889450000000,-0.027918208133030944000000,0.211190693947099300000000,0.027340263752781480000000,-0.132388305563687660000000,-0.006239722752369098900000,0.075924236044333640000000,-0.007588974368841774000000,-0.036888397691750965000000,0.010297659640913849000000,0.013993768859792647000000,-0.006990014563432881200000,-0.003644279621506338400000,0.003128023381203260100000,0.000407896980849087590000,-0.000941021749359573200000,0.000114241520038639420000,0.000174787245225280790000,-0.000061035966214111162000,-0.000013945668988208811000,0.000011336608661274467000,-0.000001043571342311495000,-0.000000736365678545024900,0.000000230878408685722150,-0.000000021093396301004384};
localparam real pDB16_Hi_D [32] = '{-0.003189220925347287500000,0.034907714323668397000000,-0.165064283488829620000000,0.430312722845942080000000,-0.637356332083695460000000,0.440290256886286200000000,0.089751089402492351000000,-0.327063310527889450000000,0.027918208133030944000000,0.211190693947099300000000,-0.027340263752781480000000,-0.132388305563687660000000,0.006239722752369098900000,0.075924236044333640000000,0.007588974368841774000000,-0.036888397691750965000000,-0.010297659640913849000000,0.013993768859792647000000,0.006990014563432881200000,-0.003644279621506338400000,-0.003128023381203260100000,0.000407896980849087590000,0.000941021749359573200000,0.000114241520038639420000,-0.000174787245225280790000,-0.000061035966214111162000,0.000013945668988208811000,0.000011336608661274467000,0.000001043571342311495000,-0.000000736365678545024900,-0.000000230878408685722150,-0.000000021093396301004384};
localparam real pDB16_Hi_R [32] = '{-0.000000021093396301004384,-0.000000230878408685722150,-0.000000736365678545024900,0.000001043571342311495000,0.000011336608661274467000,0.000013945668988208811000,-0.000061035966214111162000,-0.000174787245225280790000,0.000114241520038639420000,0.000941021749359573200000,0.000407896980849087590000,-0.003128023381203260100000,-0.003644279621506338400000,0.006990014563432881200000,0.013993768859792647000000,-0.010297659640913849000000,-0.036888397691750965000000,0.007588974368841774000000,0.075924236044333640000000,0.006239722752369098900000,-0.132388305563687660000000,-0.027340263752781480000000,0.211190693947099300000000,0.027918208133030944000000,-0.327063310527889450000000,0.089751089402492351000000,0.440290256886286200000000,-0.637356332083695460000000,0.430312722845942080000000,-0.165064283488829620000000,0.034907714323668397000000,-0.003189220925347287500000};

localparam real pDB17_Lo_D [34] = '{0.000000007267492968546472,-0.000000084239484459851937,0.000000295770093331070850,0.000000301654960998839990,-0.000004505942477213676900,0.000006990600985061646300,0.000023186813798695686000,-0.000082048032024368832000,-0.000025610109566488664000,0.000439465427767898570000,-0.000328132519408249340000,-0.001436845304796914700000,0.002301205242156734500000,0.002967996691536946700000,-0.008602921520273280500000,-0.003042989981291581700000,0.022733676584004769000000,-0.003270955535616020600000,-0.046922438388842892000000,0.022312336178527254000000,0.081105986654549503000000,-0.057091419631021115000000,-0.126815691777618340000000,0.101135489177482070000000,0.197310589564678370000000,-0.126599752215611430000000,-0.328320748363291780000000,0.027314970403216999000000,0.518315764055837790000000,0.610996615683334960000000,0.370350724151862150000000,0.131214903307548670000000,0.025985393703551473000000,0.002241807001032606900000};
localparam real pDB17_Lo_R [34] = '{0.002241807001032606900000,0.025985393703551473000000,0.131214903307548670000000,0.370350724151862150000000,0.610996615683334960000000,0.518315764055837790000000,0.027314970403216999000000,-0.328320748363291780000000,-0.126599752215611430000000,0.197310589564678370000000,0.101135489177482070000000,-0.126815691777618340000000,-0.057091419631021115000000,0.081105986654549503000000,0.022312336178527254000000,-0.046922438388842892000000,-0.003270955535616020600000,0.022733676584004769000000,-0.003042989981291581700000,-0.008602921520273280500000,0.002967996691536946700000,0.002301205242156734500000,-0.001436845304796914700000,-0.000328132519408249340000,0.000439465427767898570000,-0.000025610109566488664000,-0.000082048032024368832000,0.000023186813798695686000,0.000006990600985061646300,-0.000004505942477213676900,0.000000301654960998839990,0.000000295770093331070850,-0.000000084239484459851937,0.000000007267492968546472};
localparam real pDB17_Hi_D [34] = '{-0.002241807001032606900000,0.025985393703551473000000,-0.131214903307548670000000,0.370350724151862150000000,-0.610996615683334960000000,0.518315764055837790000000,-0.027314970403216999000000,-0.328320748363291780000000,0.126599752215611430000000,0.197310589564678370000000,-0.101135489177482070000000,-0.126815691777618340000000,0.057091419631021115000000,0.081105986654549503000000,-0.022312336178527254000000,-0.046922438388842892000000,0.003270955535616020600000,0.022733676584004769000000,0.003042989981291581700000,-0.008602921520273280500000,-0.002967996691536946700000,0.002301205242156734500000,0.001436845304796914700000,-0.000328132519408249340000,-0.000439465427767898570000,-0.000025610109566488664000,0.000082048032024368832000,0.000023186813798695686000,-0.000006990600985061646300,-0.000004505942477213676900,-0.000000301654960998839990,0.000000295770093331070850,0.000000084239484459851937,0.000000007267492968546472};
localparam real pDB17_Hi_R [34] = '{0.000000007267492968546472,0.000000084239484459851937,0.000000295770093331070850,-0.000000301654960998839990,-0.000004505942477213676900,-0.000006990600985061646300,0.000023186813798695686000,0.000082048032024368832000,-0.000025610109566488664000,-0.000439465427767898570000,-0.000328132519408249340000,0.001436845304796914700000,0.002301205242156734500000,-0.002967996691536946700000,-0.008602921520273280500000,0.003042989981291581700000,0.022733676584004769000000,0.003270955535616020600000,-0.046922438388842892000000,-0.022312336178527254000000,0.081105986654549503000000,0.057091419631021115000000,-0.126815691777618340000000,-0.101135489177482070000000,0.197310589564678370000000,0.126599752215611430000000,-0.328320748363291780000000,-0.027314970403216999000000,0.518315764055837790000000,-0.610996615683334960000000,0.370350724151862150000000,-0.131214903307548670000000,0.025985393703551473000000,-0.002241807001032606900000};

localparam real pDB18_Lo_D [36] = '{-0.000000002507934454954369,0.000000030688358630522225,-0.000000117609876703093410,-0.000000076916326899038775,0.000001768712983631628700,-0.000003332634478893568100,-0.000008520602537466953600,0.000037412378807482344000,-0.000000153591712350377960,-0.000198648552312045600000,0.000213581561911882650000,0.000628465682970796380000,-0.001340596298327426000000,-0.001118732666971648600000,0.004943343605508811700000,0.000118630033872352580000,-0.013051480946692576000000,0.006262167954147145700000,0.026670705926199838000000,-0.023733210396389887000000,-0.044526141903629801000000,0.057051247738151248000000,0.064887216211639606000000,-0.106752246660366590000000,-0.092331884151252194000000,0.167081312763510320000000,0.149533975565628220000000,-0.216480934005704260000000,-0.293654040737270030000000,0.147223111970251510000000,0.571801654889962150000000,0.571826807767921830000000,0.314678941337755590000000,0.103588465822661920000000,0.019288531724190750000000,0.001576310218444387000000};
localparam real pDB18_Lo_R [36] = '{0.001576310218444387000000,0.019288531724190750000000,0.103588465822661920000000,0.314678941337755590000000,0.571826807767921830000000,0.571801654889962150000000,0.147223111970251510000000,-0.293654040737270030000000,-0.216480934005704260000000,0.149533975565628220000000,0.167081312763510320000000,-0.092331884151252194000000,-0.106752246660366590000000,0.064887216211639606000000,0.057051247738151248000000,-0.044526141903629801000000,-0.023733210396389887000000,0.026670705926199838000000,0.006262167954147145700000,-0.013051480946692576000000,0.000118630033872352580000,0.004943343605508811700000,-0.001118732666971648600000,-0.001340596298327426000000,0.000628465682970796380000,0.000213581561911882650000,-0.000198648552312045600000,-0.000000153591712350377960,0.000037412378807482344000,-0.000008520602537466953600,-0.000003332634478893568100,0.000001768712983631628700,-0.000000076916326899038775,-0.000000117609876703093410,0.000000030688358630522225,-0.000000002507934454954369};
localparam real pDB18_Hi_D [36] = '{-0.001576310218444387000000,0.019288531724190750000000,-0.103588465822661920000000,0.314678941337755590000000,-0.571826807767921830000000,0.571801654889962150000000,-0.147223111970251510000000,-0.293654040737270030000000,0.216480934005704260000000,0.149533975565628220000000,-0.167081312763510320000000,-0.092331884151252194000000,0.106752246660366590000000,0.064887216211639606000000,-0.057051247738151248000000,-0.044526141903629801000000,0.023733210396389887000000,0.026670705926199838000000,-0.006262167954147145700000,-0.013051480946692576000000,-0.000118630033872352580000,0.004943343605508811700000,0.001118732666971648600000,-0.001340596298327426000000,-0.000628465682970796380000,0.000213581561911882650000,0.000198648552312045600000,-0.000000153591712350377960,-0.000037412378807482344000,-0.000008520602537466953600,0.000003332634478893568100,0.000001768712983631628700,0.000000076916326899038775,-0.000000117609876703093410,-0.000000030688358630522225,-0.000000002507934454954369};
localparam real pDB18_Hi_R [36] = '{-0.000000002507934454954369,-0.000000030688358630522225,-0.000000117609876703093410,0.000000076916326899038775,0.000001768712983631628700,0.000003332634478893568100,-0.000008520602537466953600,-0.000037412378807482344000,-0.000000153591712350377960,0.000198648552312045600000,0.000213581561911882650000,-0.000628465682970796380000,-0.001340596298327426000000,0.001118732666971648600000,0.004943343605508811700000,-0.000118630033872352580000,-0.013051480946692576000000,-0.006262167954147145700000,0.026670705926199838000000,0.023733210396389887000000,-0.044526141903629801000000,-0.057051247738151248000000,0.064887216211639606000000,0.106752246660366590000000,-0.092331884151252194000000,-0.167081312763510320000000,0.149533975565628220000000,0.216480934005704260000000,-0.293654040737270030000000,-0.147223111970251510000000,0.571801654889962150000000,-0.571826807767921830000000,0.314678941337755590000000,-0.103588465822661920000000,0.019288531724190750000000,-0.001576310218444387000000};

localparam real pDB19_Lo_D [38] = '{0.000000000866684883899211,-0.000000011164020670351114,0.000000046369377757796068,0.000000014470882987968016,-0.000000686275565776468310,0.000001531931476690311900,0.000003010964316295239900,-0.000016640176297141985000,0.000005105950487072856200,0.000087112704672122563000,-0.000124600791734198870000,-0.000260676135678783690000,0.000735802520504504000000,0.000341808653458229510000,-0.002687551800699482700000,0.000768954359255526010000,0.007040747367089613900000,-0.005866922281039202400000,-0.013988388678576900000000,0.019375549889116422000000,0.021623767409572607000000,-0.045674226277109146000000,-0.026501236249915492000000,0.086906755556003745000000,0.027584350625845820000000,-0.142785695038478520000000,-0.033518541902197767000000,0.212349743306165540000000,0.074652269708052124000000,-0.285838631755648550000000,-0.228091394215335530000000,0.260894952650877090000000,0.601704549127157980000000,0.524436377464322260000000,0.264388431740728740000000,0.081278113265407820000000,0.014281098450755304000000,0.001108669763181004300000};
localparam real pDB19_Lo_R [38] = '{0.001108669763181004300000,0.014281098450755304000000,0.081278113265407820000000,0.264388431740728740000000,0.524436377464322260000000,0.601704549127157980000000,0.260894952650877090000000,-0.228091394215335530000000,-0.285838631755648550000000,0.074652269708052124000000,0.212349743306165540000000,-0.033518541902197767000000,-0.142785695038478520000000,0.027584350625845820000000,0.086906755556003745000000,-0.026501236249915492000000,-0.045674226277109146000000,0.021623767409572607000000,0.019375549889116422000000,-0.013988388678576900000000,-0.005866922281039202400000,0.007040747367089613900000,0.000768954359255526010000,-0.002687551800699482700000,0.000341808653458229510000,0.000735802520504504000000,-0.000260676135678783690000,-0.000124600791734198870000,0.000087112704672122563000,0.000005105950487072856200,-0.000016640176297141985000,0.000003010964316295239900,0.000001531931476690311900,-0.000000686275565776468310,0.000000014470882987968016,0.000000046369377757796068,-0.000000011164020670351114,0.000000000866684883899211};
localparam real pDB19_Hi_D [38] = '{-0.001108669763181004300000,0.014281098450755304000000,-0.081278113265407820000000,0.264388431740728740000000,-0.524436377464322260000000,0.601704549127157980000000,-0.260894952650877090000000,-0.228091394215335530000000,0.285838631755648550000000,0.074652269708052124000000,-0.212349743306165540000000,-0.033518541902197767000000,0.142785695038478520000000,0.027584350625845820000000,-0.086906755556003745000000,-0.026501236249915492000000,0.045674226277109146000000,0.021623767409572607000000,-0.019375549889116422000000,-0.013988388678576900000000,0.005866922281039202400000,0.007040747367089613900000,-0.000768954359255526010000,-0.002687551800699482700000,-0.000341808653458229510000,0.000735802520504504000000,0.000260676135678783690000,-0.000124600791734198870000,-0.000087112704672122563000,0.000005105950487072856200,0.000016640176297141985000,0.000003010964316295239900,-0.000001531931476690311900,-0.000000686275565776468310,-0.000000014470882987968016,0.000000046369377757796068,0.000000011164020670351114,0.000000000866684883899211};
localparam real pDB19_Hi_R [38] = '{0.000000000866684883899211,0.000000011164020670351114,0.000000046369377757796068,-0.000000014470882987968016,-0.000000686275565776468310,-0.000001531931476690311900,0.000003010964316295239900,0.000016640176297141985000,0.000005105950487072856200,-0.000087112704672122563000,-0.000124600791734198870000,0.000260676135678783690000,0.000735802520504504000000,-0.000341808653458229510000,-0.002687551800699482700000,-0.000768954359255526010000,0.007040747367089613900000,0.005866922281039202400000,-0.013988388678576900000000,-0.019375549889116422000000,0.021623767409572607000000,0.045674226277109146000000,-0.026501236249915492000000,-0.086906755556003745000000,0.027584350625845820000000,0.142785695038478520000000,-0.033518541902197767000000,-0.212349743306165540000000,0.074652269708052124000000,0.285838631755648550000000,-0.228091394215335530000000,-0.260894952650877090000000,0.601704549127157980000000,-0.524436377464322260000000,0.264388431740728740000000,-0.081278113265407820000000,0.014281098450755304000000,-0.001108669763181004300000};

localparam real pDB20_Lo_D [40] = '{-0.000000000299883648961136,0.000000004056127055541042,-0.000000018148432482948567,0.000000000201432202355199,0.000000263392422626301800,-0.000000684707959698251880,-0.000001011994010016522700,0.000007241248287651389200,-0.000004376143862191575500,-0.000037105861833940264000,0.000067742808283264108000,0.000101532889735460870000,-0.000385104748700683310000,-0.000053497598446011665000,0.001392559619303886600000,-0.000831562172857963940000,-0.003581494259679262200000,0.004420542386902407200000,0.006721627302091013600000,-0.013810526137172797000000,-0.008789324923671099100000,0.032294299531286479000000,0.005874681812756509300000,-0.061722899623438486000000,0.005632246858176481700000,0.102291719174675010000000,-0.024716827338396870000000,-0.155458750706898990000000,0.039850246457581083000000,0.228291050819266320000000,-0.016727088309026167000000,-0.326786800433140120000000,-0.139212088011097380000000,0.361502298738368920000000,0.610493238936961390000000,0.472696185309637200000000,0.219942113550808750000000,0.063423780458911894000000,0.010549394624922191000000,0.000779953613664761260000};
localparam real pDB20_Lo_R [40] = '{0.000779953613664761260000,0.010549394624922191000000,0.063423780458911894000000,0.219942113550808750000000,0.472696185309637200000000,0.610493238936961390000000,0.361502298738368920000000,-0.139212088011097380000000,-0.326786800433140120000000,-0.016727088309026167000000,0.228291050819266320000000,0.039850246457581083000000,-0.155458750706898990000000,-0.024716827338396870000000,0.102291719174675010000000,0.005632246858176481700000,-0.061722899623438486000000,0.005874681812756509300000,0.032294299531286479000000,-0.008789324923671099100000,-0.013810526137172797000000,0.006721627302091013600000,0.004420542386902407200000,-0.003581494259679262200000,-0.000831562172857963940000,0.001392559619303886600000,-0.000053497598446011665000,-0.000385104748700683310000,0.000101532889735460870000,0.000067742808283264108000,-0.000037105861833940264000,-0.000004376143862191575500,0.000007241248287651389200,-0.000001011994010016522700,-0.000000684707959698251880,0.000000263392422626301800,0.000000000201432202355199,-0.000000018148432482948567,0.000000004056127055541042,-0.000000000299883648961136};
localparam real pDB20_Hi_D [40] = '{-0.000779953613664761260000,0.010549394624922191000000,-0.063423780458911894000000,0.219942113550808750000000,-0.472696185309637200000000,0.610493238936961390000000,-0.361502298738368920000000,-0.139212088011097380000000,0.326786800433140120000000,-0.016727088309026167000000,-0.228291050819266320000000,0.039850246457581083000000,0.155458750706898990000000,-0.024716827338396870000000,-0.102291719174675010000000,0.005632246858176481700000,0.061722899623438486000000,0.005874681812756509300000,-0.032294299531286479000000,-0.008789324923671099100000,0.013810526137172797000000,0.006721627302091013600000,-0.004420542386902407200000,-0.003581494259679262200000,0.000831562172857963940000,0.001392559619303886600000,0.000053497598446011665000,-0.000385104748700683310000,-0.000101532889735460870000,0.000067742808283264108000,0.000037105861833940264000,-0.000004376143862191575500,-0.000007241248287651389200,-0.000001011994010016522700,0.000000684707959698251880,0.000000263392422626301800,-0.000000000201432202355199,-0.000000018148432482948567,-0.000000004056127055541042,-0.000000000299883648961136};
localparam real pDB20_Hi_R [40] = '{-0.000000000299883648961136,-0.000000004056127055541042,-0.000000018148432482948567,-0.000000000201432202355199,0.000000263392422626301800,0.000000684707959698251880,-0.000001011994010016522700,-0.000007241248287651389200,-0.000004376143862191575500,0.000037105861833940264000,0.000067742808283264108000,-0.000101532889735460870000,-0.000385104748700683310000,0.000053497598446011665000,0.001392559619303886600000,0.000831562172857963940000,-0.003581494259679262200000,-0.004420542386902407200000,0.006721627302091013600000,0.013810526137172797000000,-0.008789324923671099100000,-0.032294299531286479000000,0.005874681812756509300000,0.061722899623438486000000,0.005632246858176481700000,-0.102291719174675010000000,-0.024716827338396870000000,0.155458750706898990000000,0.039850246457581083000000,-0.228291050819266320000000,-0.016727088309026167000000,0.326786800433140120000000,-0.139212088011097380000000,-0.361502298738368920000000,0.610493238936961390000000,-0.472696185309637200000000,0.219942113550808750000000,-0.063423780458911894000000,0.010549394624922191000000,-0.000779953613664761260000};

localparam real pCOIF1_Lo_D [6] = '{-0.015655728135464540000000,-0.072732619512853897000000,0.384864846864202860000000,0.852572020212255420000000,0.337897662457809220000000,-0.072732619512853897000000};
localparam real pCOIF1_Lo_R [6] = '{-0.072732619512853897000000,0.337897662457809220000000,0.852572020212255420000000,0.384864846864202860000000,-0.072732619512853897000000,-0.015655728135464540000000};
localparam real pCOIF1_Hi_D [6] = '{0.072732619512853897000000,0.337897662457809220000000,-0.852572020212255420000000,0.384864846864202860000000,0.072732619512853897000000,-0.015655728135464540000000};
localparam real pCOIF1_Hi_R [6] = '{-0.015655728135464540000000,0.072732619512853897000000,0.384864846864202860000000,-0.852572020212255420000000,0.337897662457809220000000,0.072732619512853897000000};

localparam real pCOIF2_Lo_D [12] = '{-0.000720549445364512210000,-0.001823208870702993200000,0.005611434819394499500000,0.023680171946334084000000,-0.059434418646456898000000,-0.076488599078306393000000,0.417005184421692540000000,0.812723635445542270000000,0.386110066821162220000000,-0.067372554721963018000000,-0.041464936781759151000000,0.016387336463522112000000};
localparam real pCOIF2_Lo_R [12] = '{0.016387336463522112000000,-0.041464936781759151000000,-0.067372554721963018000000,0.386110066821162220000000,0.812723635445542270000000,0.417005184421692540000000,-0.076488599078306393000000,-0.059434418646456898000000,0.023680171946334084000000,0.005611434819394499500000,-0.001823208870702993200000,-0.000720549445364512210000};
localparam real pCOIF2_Hi_D [12] = '{-0.016387336463522112000000,-0.041464936781759151000000,0.067372554721963018000000,0.386110066821162220000000,-0.812723635445542270000000,0.417005184421692540000000,0.076488599078306393000000,-0.059434418646456898000000,-0.023680171946334084000000,0.005611434819394499500000,0.001823208870702993200000,-0.000720549445364512210000};
localparam real pCOIF2_Hi_R [12] = '{-0.000720549445364512210000,0.001823208870702993200000,0.005611434819394499500000,-0.023680171946334084000000,-0.059434418646456898000000,0.076488599078306393000000,0.417005184421692540000000,-0.812723635445542270000000,0.386110066821162220000000,0.067372554721963018000000,-0.041464936781759151000000,-0.016387336463522112000000};

localparam real pCOIF3_Lo_D [18] = '{-0.000034599772836212559000,-0.000070983303138141252000,0.000466216960112886310000,0.001117518770890601600000,-0.002574517688750223600000,-0.009007976136661580500000,0.015880544863615904000000,0.034555027573061628000000,-0.082301927106885983000000,-0.071799821619312018000000,0.428483476377618740000000,0.793777222625620560000000,0.405176902409616900000000,-0.061123390002672869000000,-0.065771911281855500000000,0.023452696141836267000000,0.007782596427325418200000,-0.003793512864491014100000};
localparam real pCOIF3_Lo_R [18] = '{-0.003793512864491014100000,0.007782596427325418200000,0.023452696141836267000000,-0.065771911281855500000000,-0.061123390002672869000000,0.405176902409616900000000,0.793777222625620560000000,0.428483476377618740000000,-0.071799821619312018000000,-0.082301927106885983000000,0.034555027573061628000000,0.015880544863615904000000,-0.009007976136661580500000,-0.002574517688750223600000,0.001117518770890601600000,0.000466216960112886310000,-0.000070983303138141252000,-0.000034599772836212559000};
localparam real pCOIF3_Hi_D [18] = '{0.003793512864491014100000,0.007782596427325418200000,-0.023452696141836267000000,-0.065771911281855500000000,0.061123390002672869000000,0.405176902409616900000000,-0.793777222625620560000000,0.428483476377618740000000,0.071799821619312018000000,-0.082301927106885983000000,-0.034555027573061628000000,0.015880544863615904000000,0.009007976136661580500000,-0.002574517688750223600000,-0.001117518770890601600000,0.000466216960112886310000,0.000070983303138141252000,-0.000034599772836212559000};
localparam real pCOIF3_Hi_R [18] = '{-0.000034599772836212559000,0.000070983303138141252000,0.000466216960112886310000,-0.001117518770890601600000,-0.002574517688750223600000,0.009007976136661580500000,0.015880544863615904000000,-0.034555027573061628000000,-0.082301927106885983000000,0.071799821619312018000000,0.428483476377618740000000,-0.793777222625620560000000,0.405176902409616900000000,0.061123390002672869000000,-0.065771911281855500000000,-0.023452696141836267000000,0.007782596427325418200000,0.003793512864491014100000};

localparam real pCOIF4_Lo_D [24] = '{-0.000001784985003088261400,-0.000003259680236883367500,0.000031229875865345646000,0.000062339034461007128000,-0.000259974552487713240000,-0.000589020756244338310000,0.001266561929298944500000,0.003751436157278457100000,-0.005658286686610719900000,-0.015211731527946259000000,0.025082261844864097000000,0.039334427123337491000000,-0.096220442033987982000000,-0.066627474263425038000000,0.434386056491468500000000,0.782238930920499010000000,0.415308407030430260000000,-0.056077313316754807000000,-0.081266699680878754000000,0.026682300156053072000000,0.016068943964776348000000,-0.007346166327642093500000,-0.001629492012601732600000,0.000892313668582314560000};
localparam real pCOIF4_Lo_R [24] = '{0.000892313668582314560000,-0.001629492012601732600000,-0.007346166327642093500000,0.016068943964776348000000,0.026682300156053072000000,-0.081266699680878754000000,-0.056077313316754807000000,0.415308407030430260000000,0.782238930920499010000000,0.434386056491468500000000,-0.066627474263425038000000,-0.096220442033987982000000,0.039334427123337491000000,0.025082261844864097000000,-0.015211731527946259000000,-0.005658286686610719900000,0.003751436157278457100000,0.001266561929298944500000,-0.000589020756244338310000,-0.000259974552487713240000,0.000062339034461007128000,0.000031229875865345646000,-0.000003259680236883367500,-0.000001784985003088261400};
localparam real pCOIF4_Hi_D [24] = '{-0.000892313668582314560000,-0.001629492012601732600000,0.007346166327642093500000,0.016068943964776348000000,-0.026682300156053072000000,-0.081266699680878754000000,0.056077313316754807000000,0.415308407030430260000000,-0.782238930920499010000000,0.434386056491468500000000,0.066627474263425038000000,-0.096220442033987982000000,-0.039334427123337491000000,0.025082261844864097000000,0.015211731527946259000000,-0.005658286686610719900000,-0.003751436157278457100000,0.001266561929298944500000,0.000589020756244338310000,-0.000259974552487713240000,-0.000062339034461007128000,0.000031229875865345646000,0.000003259680236883367500,-0.000001784985003088261400};
localparam real pCOIF4_Hi_R [24] = '{-0.000001784985003088261400,0.000003259680236883367500,0.000031229875865345646000,-0.000062339034461007128000,-0.000259974552487713240000,0.000589020756244338310000,0.001266561929298944500000,-0.003751436157278457100000,-0.005658286686610719900000,0.015211731527946259000000,0.025082261844864097000000,-0.039334427123337491000000,-0.096220442033987982000000,0.066627474263425038000000,0.434386056491468500000000,-0.782238930920499010000000,0.415308407030430260000000,0.056077313316754807000000,-0.081266699680878754000000,-0.026682300156053072000000,0.016068943964776348000000,0.007346166327642093500000,-0.001629492012601732600000,-0.000892313668582314560000};

localparam real pCOIF5_Lo_D [30] = '{-0.000000095176572738191650,-0.000000167442885768230170,0.000002063761851364681400,0.000003734655175141404700,-0.000021315026809955787000,-0.000041340432272512511000,0.000140541149702034370000,0.000302259581813063150000,-0.000638131343045111420000,-0.001662863702013083800000,0.002433373212657672200000,0.006764185448053083200000,-0.009164231162481845800000,-0.019761778942572639000000,0.032683574267111833000000,0.041289208750181702000000,-0.105574208703338930000000,-0.062035963962903569000000,0.437991626171837120000000,0.774289603652956180000000,0.421566206690851490000000,-0.052043163176243773000000,-0.091920010559696244000000,0.028168028970936350000000,0.023408156785839195000000,-0.010131117519849788000000,-0.004159358781386048000000,0.002178236358109017800000,0.000358589687895737850000,-0.000212080839803798270000};
localparam real pCOIF5_Lo_R [30] = '{-0.000212080839803798270000,0.000358589687895737850000,0.002178236358109017800000,-0.004159358781386048000000,-0.010131117519849788000000,0.023408156785839195000000,0.028168028970936350000000,-0.091920010559696244000000,-0.052043163176243773000000,0.421566206690851490000000,0.774289603652956180000000,0.437991626171837120000000,-0.062035963962903569000000,-0.105574208703338930000000,0.041289208750181702000000,0.032683574267111833000000,-0.019761778942572639000000,-0.009164231162481845800000,0.006764185448053083200000,0.002433373212657672200000,-0.001662863702013083800000,-0.000638131343045111420000,0.000302259581813063150000,0.000140541149702034370000,-0.000041340432272512511000,-0.000021315026809955787000,0.000003734655175141404700,0.000002063761851364681400,-0.000000167442885768230170,-0.000000095176572738191650};
localparam real pCOIF5_Hi_D [30] = '{0.000212080839803798270000,0.000358589687895737850000,-0.002178236358109017800000,-0.004159358781386048000000,0.010131117519849788000000,0.023408156785839195000000,-0.028168028970936350000000,-0.091920010559696244000000,0.052043163176243773000000,0.421566206690851490000000,-0.774289603652956180000000,0.437991626171837120000000,0.062035963962903569000000,-0.105574208703338930000000,-0.041289208750181702000000,0.032683574267111833000000,0.019761778942572639000000,-0.009164231162481845800000,-0.006764185448053083200000,0.002433373212657672200000,0.001662863702013083800000,-0.000638131343045111420000,-0.000302259581813063150000,0.000140541149702034370000,0.000041340432272512511000,-0.000021315026809955787000,-0.000003734655175141404700,0.000002063761851364681400,0.000000167442885768230170,-0.000000095176572738191650};
localparam real pCOIF5_Hi_R [30] = '{-0.000000095176572738191650,0.000000167442885768230170,0.000002063761851364681400,-0.000003734655175141404700,-0.000021315026809955787000,0.000041340432272512511000,0.000140541149702034370000,-0.000302259581813063150000,-0.000638131343045111420000,0.001662863702013083800000,0.002433373212657672200000,-0.006764185448053083200000,-0.009164231162481845800000,0.019761778942572639000000,0.032683574267111833000000,-0.041289208750181702000000,-0.105574208703338930000000,0.062035963962903569000000,0.437991626171837120000000,-0.774289603652956180000000,0.421566206690851490000000,0.052043163176243773000000,-0.091920010559696244000000,-0.028168028970936350000000,0.023408156785839195000000,0.010131117519849788000000,-0.004159358781386048000000,-0.002178236358109017800000,0.000358589687895737850000,0.000212080839803798270000};

localparam real pSYM2_Lo_D [4] = '{-0.129409522550921450000000,0.224143868041857350000000,0.836516303737468990000000,0.482962913144690250000000};
localparam real pSYM2_Lo_R [4] = '{0.482962913144690250000000,0.836516303737468990000000,0.224143868041857350000000,-0.129409522550921450000000};
localparam real pSYM2_Hi_D [4] = '{-0.482962913144690250000000,0.836516303737468990000000,-0.224143868041857350000000,-0.129409522550921450000000};
localparam real pSYM2_Hi_R [4] = '{-0.129409522550921450000000,-0.224143868041857350000000,0.836516303737468990000000,-0.482962913144690250000000};

localparam real pSYM3_Lo_D [6] = '{0.035226291882100656000000,-0.085441273882241486000000,-0.135011020010390840000000,0.459877502119331320000000,0.806891509313338750000000,0.332670552950956880000000};
localparam real pSYM3_Lo_R [6] = '{0.332670552950956880000000,0.806891509313338750000000,0.459877502119331320000000,-0.135011020010390840000000,-0.085441273882241486000000,0.035226291882100656000000};
localparam real pSYM3_Hi_D [6] = '{-0.332670552950956880000000,0.806891509313338750000000,-0.459877502119331320000000,-0.135011020010390840000000,0.085441273882241486000000,0.035226291882100656000000};
localparam real pSYM3_Hi_R [6] = '{0.035226291882100656000000,0.085441273882241486000000,-0.135011020010390840000000,-0.459877502119331320000000,0.806891509313338750000000,-0.332670552950956880000000};

localparam real pSYM4_Lo_D [8] = '{-0.075765714789273325000000,-0.029635527645998510000000,0.497618667632015450000000,0.803738751805916140000000,0.297857795605277360000000,-0.099219543576847216000000,-0.012603967262037833000000,0.032223100604042702000000};
localparam real pSYM4_Lo_R [8] = '{0.032223100604042702000000,-0.012603967262037833000000,-0.099219543576847216000000,0.297857795605277360000000,0.803738751805916140000000,0.497618667632015450000000,-0.029635527645998510000000,-0.075765714789273325000000};
localparam real pSYM4_Hi_D [8] = '{-0.032223100604042702000000,-0.012603967262037833000000,0.099219543576847216000000,0.297857795605277360000000,-0.803738751805916140000000,0.497618667632015450000000,0.029635527645998510000000,-0.075765714789273325000000};
localparam real pSYM4_Hi_R [8] = '{-0.075765714789273325000000,0.029635527645998510000000,0.497618667632015450000000,-0.803738751805916140000000,0.297857795605277360000000,0.099219543576847216000000,-0.012603967262037833000000,-0.032223100604042702000000};

localparam real pSYM5_Lo_D [10] = '{0.027333068345077982000000,0.029519490925774643000000,-0.039134249302383094000000,0.199397533977393600000000,0.723407690402420590000000,0.633978963458211920000000,0.016602105764522319000000,-0.175328089908450470000000,-0.021101834024758855000000,0.019538882735286728000000};
localparam real pSYM5_Lo_R [10] = '{0.019538882735286728000000,-0.021101834024758855000000,-0.175328089908450470000000,0.016602105764522319000000,0.633978963458211920000000,0.723407690402420590000000,0.199397533977393600000000,-0.039134249302383094000000,0.029519490925774643000000,0.027333068345077982000000};
localparam real pSYM5_Hi_D [10] = '{-0.019538882735286728000000,-0.021101834024758855000000,0.175328089908450470000000,0.016602105764522319000000,-0.633978963458211920000000,0.723407690402420590000000,-0.199397533977393600000000,-0.039134249302383094000000,-0.029519490925774643000000,0.027333068345077982000000};
localparam real pSYM5_Hi_R [10] = '{0.027333068345077982000000,-0.029519490925774643000000,-0.039134249302383094000000,-0.199397533977393600000000,0.723407690402420590000000,-0.633978963458211920000000,0.016602105764522319000000,0.175328089908450470000000,-0.021101834024758855000000,-0.019538882735286728000000};

localparam real pSYM6_Lo_D [12] = '{0.015404109327027373000000,0.003490712084217470200000,-0.117990111148190570000000,-0.048311742585632998000000,0.491055941926746620000000,0.787641141030194000000000,0.337929421727621800000000,-0.072637522786462516000000,-0.021060292512300564000000,0.044724901770665779000000,0.001767711864242803600000,-0.007800708325034148000000};
localparam real pSYM6_Lo_R [12] = '{-0.007800708325034148000000,0.001767711864242803600000,0.044724901770665779000000,-0.021060292512300564000000,-0.072637522786462516000000,0.337929421727621800000000,0.787641141030194000000000,0.491055941926746620000000,-0.048311742585632998000000,-0.117990111148190570000000,0.003490712084217470200000,0.015404109327027373000000};
localparam real pSYM6_Hi_D [12] = '{0.007800708325034148000000,0.001767711864242803600000,-0.044724901770665779000000,-0.021060292512300564000000,0.072637522786462516000000,0.337929421727621800000000,-0.787641141030194000000000,0.491055941926746620000000,0.048311742585632998000000,-0.117990111148190570000000,-0.003490712084217470200000,0.015404109327027373000000};
localparam real pSYM6_Hi_R [12] = '{0.015404109327027373000000,-0.003490712084217470200000,-0.117990111148190570000000,0.048311742585632998000000,0.491055941926746620000000,-0.787641141030194000000000,0.337929421727621800000000,0.072637522786462516000000,-0.021060292512300564000000,-0.044724901770665779000000,0.001767711864242803600000,0.007800708325034148000000};

localparam real pSYM7_Lo_D [14] = '{0.002681814568257878100000,-0.001047384888682916300000,-0.012636303403251930000000,0.030515513165963570000000,0.067892693501372697000000,-0.049552834937127255000000,0.017441255086855827000000,0.536101917091762800000000,0.767764317003164050000000,0.288629631751514630000000,-0.140047240442961520000000,-0.107808237703817740000000,0.004010244871533663400000,0.010268176708511255000000};
localparam real pSYM7_Lo_R [14] = '{0.010268176708511255000000,0.004010244871533663400000,-0.107808237703817740000000,-0.140047240442961520000000,0.288629631751514630000000,0.767764317003164050000000,0.536101917091762800000000,0.017441255086855827000000,-0.049552834937127255000000,0.067892693501372697000000,0.030515513165963570000000,-0.012636303403251930000000,-0.001047384888682916300000,0.002681814568257878100000};
localparam real pSYM7_Hi_D [14] = '{-0.010268176708511255000000,0.004010244871533663400000,0.107808237703817740000000,-0.140047240442961520000000,-0.288629631751514630000000,0.767764317003164050000000,-0.536101917091762800000000,0.017441255086855827000000,0.049552834937127255000000,0.067892693501372697000000,-0.030515513165963570000000,-0.012636303403251930000000,0.001047384888682916300000,0.002681814568257878100000};
localparam real pSYM7_Hi_R [14] = '{0.002681814568257878100000,0.001047384888682916300000,-0.012636303403251930000000,-0.030515513165963570000000,0.067892693501372697000000,0.049552834937127255000000,0.017441255086855827000000,-0.536101917091762800000000,0.767764317003164050000000,-0.288629631751514630000000,-0.140047240442961520000000,0.107808237703817740000000,0.004010244871533663400000,-0.010268176708511255000000};

localparam real pSYM8_Lo_D [16] = '{-0.003382415951006125600000,-0.000542132331791148120000,0.031695087811492981000000,0.007607487324917605400000,-0.143294238350809710000000,-0.061273359067658524000000,0.481359651258372210000000,0.777185751700523510000000,0.364441894835331400000000,-0.051945838107709037000000,-0.027219029917056003000000,0.049137179673607506000000,0.003808752013890615100000,-0.014952258337048231000000,-0.000302920514721366800000,0.001889950332759460900000};
localparam real pSYM8_Lo_R [16] = '{0.001889950332759460900000,-0.000302920514721366800000,-0.014952258337048231000000,0.003808752013890615100000,0.049137179673607506000000,-0.027219029917056003000000,-0.051945838107709037000000,0.364441894835331400000000,0.777185751700523510000000,0.481359651258372210000000,-0.061273359067658524000000,-0.143294238350809710000000,0.007607487324917605400000,0.031695087811492981000000,-0.000542132331791148120000,-0.003382415951006125600000};
localparam real pSYM8_Hi_D [16] = '{-0.001889950332759460900000,-0.000302920514721366800000,0.014952258337048231000000,0.003808752013890615100000,-0.049137179673607506000000,-0.027219029917056003000000,0.051945838107709037000000,0.364441894835331400000000,-0.777185751700523510000000,0.481359651258372210000000,0.061273359067658524000000,-0.143294238350809710000000,-0.007607487324917605400000,0.031695087811492981000000,0.000542132331791148120000,-0.003382415951006125600000};
localparam real pSYM8_Hi_R [16] = '{-0.003382415951006125600000,0.000542132331791148120000,0.031695087811492981000000,-0.007607487324917605400000,-0.143294238350809710000000,0.061273359067658524000000,0.481359651258372210000000,-0.777185751700523510000000,0.364441894835331400000000,0.051945838107709037000000,-0.027219029917056003000000,-0.049137179673607506000000,0.003808752013890615100000,0.014952258337048231000000,-0.000302920514721366800000,-0.001889950332759460900000};

localparam real pSYM9_Lo_D [18] = '{0.001400915525914665300000,0.000619780888985553800000,-0.013271967781817105000000,-0.011528210207679338000000,0.030224878858275173000000,0.000583462746125848260000,-0.054568958430832502000000,0.238760914607303840000000,0.717897082764410110000000,0.617338449140934500000000,0.035272488035273511000000,-0.191550831297283420000000,-0.018233770779396471000000,0.062077789302885017000000,0.008859267493400243100000,-0.010264064027633073000000,-0.000473154498680074000000,0.001069490032908597500000};
localparam real pSYM9_Lo_R [18] = '{0.001069490032908597500000,-0.000473154498680074000000,-0.010264064027633073000000,0.008859267493400243100000,0.062077789302885017000000,-0.018233770779396471000000,-0.191550831297283420000000,0.035272488035273511000000,0.617338449140934500000000,0.717897082764410110000000,0.238760914607303840000000,-0.054568958430832502000000,0.000583462746125848260000,0.030224878858275173000000,-0.011528210207679338000000,-0.013271967781817105000000,0.000619780888985553800000,0.001400915525914665300000};
localparam real pSYM9_Hi_D [18] = '{-0.001069490032908597500000,-0.000473154498680074000000,0.010264064027633073000000,0.008859267493400243100000,-0.062077789302885017000000,-0.018233770779396471000000,0.191550831297283420000000,0.035272488035273511000000,-0.617338449140934500000000,0.717897082764410110000000,-0.238760914607303840000000,-0.054568958430832502000000,-0.000583462746125848260000,0.030224878858275173000000,0.011528210207679338000000,-0.013271967781817105000000,-0.000619780888985553800000,0.001400915525914665300000};
localparam real pSYM9_Hi_R [18] = '{0.001400915525914665300000,-0.000619780888985553800000,-0.013271967781817105000000,0.011528210207679338000000,0.030224878858275173000000,-0.000583462746125848260000,-0.054568958430832502000000,-0.238760914607303840000000,0.717897082764410110000000,-0.617338449140934500000000,0.035272488035273511000000,0.191550831297283420000000,-0.018233770779396471000000,-0.062077789302885017000000,0.008859267493400243100000,0.010264064027633073000000,-0.000473154498680074000000,-0.001069490032908597500000};

localparam real pSYM10_Lo_D [20] = '{0.000770159809114478620000,0.000095632670722893358000,-0.008641299277022278200000,-0.001465382581304899700000,0.045927239231092098000000,0.011609893903712620000000,-0.159494278884912880000000,-0.070880535783239690000000,0.471690666938436140000000,0.769510037021100210000000,0.383826761067083470000000,-0.035536740473815255000000,-0.031990056882427093000000,0.049994972077375743000000,0.005764912033581722100000,-0.020354939812311016000000,-0.000804358932016546970000,0.004593173585311763300000,0.000057036083618500559000,-0.000459329421004650220000};
localparam real pSYM10_Lo_R [20] = '{-0.000459329421004650220000,0.000057036083618500559000,0.004593173585311763300000,-0.000804358932016546970000,-0.020354939812311016000000,0.005764912033581722100000,0.049994972077375743000000,-0.031990056882427093000000,-0.035536740473815255000000,0.383826761067083470000000,0.769510037021100210000000,0.471690666938436140000000,-0.070880535783239690000000,-0.159494278884912880000000,0.011609893903712620000000,0.045927239231092098000000,-0.001465382581304899700000,-0.008641299277022278200000,0.000095632670722893358000,0.000770159809114478620000};
localparam real pSYM10_Hi_D [20] = '{0.000459329421004650220000,0.000057036083618500559000,-0.004593173585311763300000,-0.000804358932016546970000,0.020354939812311016000000,0.005764912033581722100000,-0.049994972077375743000000,-0.031990056882427093000000,0.035536740473815255000000,0.383826761067083470000000,-0.769510037021100210000000,0.471690666938436140000000,0.070880535783239690000000,-0.159494278884912880000000,-0.011609893903712620000000,0.045927239231092098000000,0.001465382581304899700000,-0.008641299277022278200000,-0.000095632670722893358000,0.000770159809114478620000};
localparam real pSYM10_Hi_R [20] = '{0.000770159809114478620000,-0.000095632670722893358000,-0.008641299277022278200000,0.001465382581304899700000,0.045927239231092098000000,-0.011609893903712620000000,-0.159494278884912880000000,0.070880535783239690000000,0.471690666938436140000000,-0.769510037021100210000000,0.383826761067083470000000,0.035536740473815255000000,-0.031990056882427093000000,-0.049994972077375743000000,0.005764912033581722100000,0.020354939812311016000000,-0.000804358932016546970000,-0.004593173585311763300000,0.000057036083618500559000,0.000459329421004650220000};

localparam real pSYM11_Lo_D [22] = '{0.000171721950699344420000,-0.000038795655736161771000,-0.001734366267297828000000,0.000588352735397057150000,0.006512495674771526900000,-0.009857934828789140200000,-0.024080841595862452000000,0.037037415978860080000000,0.069976799610732859000000,-0.022832651022563245000000,0.097198394458909751000000,0.572022978010083060000000,0.730343549088388060000000,0.237689909049246560000000,-0.204654794495795490000000,-0.144602343705310030000000,0.035266759564468529000000,0.043000190681552364000000,-0.002003471900109373000000,-0.006389603666454813900000,0.000110535097642741340000,0.000489263610261923120000};
localparam real pSYM11_Lo_R [22] = '{0.000489263610261923120000,0.000110535097642741340000,-0.006389603666454813900000,-0.002003471900109373000000,0.043000190681552364000000,0.035266759564468529000000,-0.144602343705310030000000,-0.204654794495795490000000,0.237689909049246560000000,0.730343549088388060000000,0.572022978010083060000000,0.097198394458909751000000,-0.022832651022563245000000,0.069976799610732859000000,0.037037415978860080000000,-0.024080841595862452000000,-0.009857934828789140200000,0.006512495674771526900000,0.000588352735397057150000,-0.001734366267297828000000,-0.000038795655736161771000,0.000171721950699344420000};
localparam real pSYM11_Hi_D [22] = '{-0.000489263610261923120000,0.000110535097642741340000,0.006389603666454813900000,-0.002003471900109373000000,-0.043000190681552364000000,0.035266759564468529000000,0.144602343705310030000000,-0.204654794495795490000000,-0.237689909049246560000000,0.730343549088388060000000,-0.572022978010083060000000,0.097198394458909751000000,0.022832651022563245000000,0.069976799610732859000000,-0.037037415978860080000000,-0.024080841595862452000000,0.009857934828789140200000,0.006512495674771526900000,-0.000588352735397057150000,-0.001734366267297828000000,0.000038795655736161771000,0.000171721950699344420000};
localparam real pSYM11_Hi_R [22] = '{0.000171721950699344420000,0.000038795655736161771000,-0.001734366267297828000000,-0.000588352735397057150000,0.006512495674771526900000,0.009857934828789140200000,-0.024080841595862452000000,-0.037037415978860080000000,0.069976799610732859000000,0.022832651022563245000000,0.097198394458909751000000,-0.572022978010083060000000,0.730343549088388060000000,-0.237689909049246560000000,-0.204654794495795490000000,0.144602343705310030000000,0.035266759564468529000000,-0.043000190681552364000000,-0.002003471900109373000000,0.006389603666454813900000,0.000110535097642741340000,-0.000489263610261923120000};

localparam real pSYM12_Lo_D [24] = '{0.000111967194246570920000,-0.000011353928041518001000,-0.001349755755571622900000,0.000180214090085178190000,0.007414965517654525900000,-0.001408909244329211900000,-0.024220722675014954000000,0.007553780611677254400000,0.049179318299659346000000,-0.035848830736960699000000,-0.022162306170360756000000,0.398885972390194130000000,0.763479097783659850000000,0.462741031219302770000000,-0.078332622316317990000000,-0.170370697238860310000000,0.015301740622475773000000,0.057804179445505602000000,-0.002604391031330956700000,-0.014589836449233978000000,0.000307647796310326520000,0.002350297614183388900000,-0.000018158078862603281000,-0.000179066586975081440000};
localparam real pSYM12_Lo_R [24] = '{-0.000179066586975081440000,-0.000018158078862603281000,0.002350297614183388900000,0.000307647796310326520000,-0.014589836449233978000000,-0.002604391031330956700000,0.057804179445505602000000,0.015301740622475773000000,-0.170370697238860310000000,-0.078332622316317990000000,0.462741031219302770000000,0.763479097783659850000000,0.398885972390194130000000,-0.022162306170360756000000,-0.035848830736960699000000,0.049179318299659346000000,0.007553780611677254400000,-0.024220722675014954000000,-0.001408909244329211900000,0.007414965517654525900000,0.000180214090085178190000,-0.001349755755571622900000,-0.000011353928041518001000,0.000111967194246570920000};
localparam real pSYM12_Hi_D [24] = '{0.000179066586975081440000,-0.000018158078862603281000,-0.002350297614183388900000,0.000307647796310326520000,0.014589836449233978000000,-0.002604391031330956700000,-0.057804179445505602000000,0.015301740622475773000000,0.170370697238860310000000,-0.078332622316317990000000,-0.462741031219302770000000,0.763479097783659850000000,-0.398885972390194130000000,-0.022162306170360756000000,0.035848830736960699000000,0.049179318299659346000000,-0.007553780611677254400000,-0.024220722675014954000000,0.001408909244329211900000,0.007414965517654525900000,-0.000180214090085178190000,-0.001349755755571622900000,0.000011353928041518001000,0.000111967194246570920000};
localparam real pSYM12_Hi_R [24] = '{0.000111967194246570920000,0.000011353928041518001000,-0.001349755755571622900000,-0.000180214090085178190000,0.007414965517654525900000,0.001408909244329211900000,-0.024220722675014954000000,-0.007553780611677254400000,0.049179318299659346000000,0.035848830736960699000000,-0.022162306170360756000000,-0.398885972390194130000000,0.763479097783659850000000,-0.462741031219302770000000,-0.078332622316317990000000,0.170370697238860310000000,0.015301740622475773000000,-0.057804179445505602000000,-0.002604391031330956700000,0.014589836449233978000000,0.000307647796310326520000,-0.002350297614183388900000,-0.000018158078862603281000,0.000179066586975081440000};

localparam real pSYM13_Lo_D [26] = '{0.000068203252630752971000,-0.000035738623648692444000,-0.001136063438928119200000,-0.000170942858530178690000,0.007526225389968108300000,0.005296359738724500500000,-0.020216768133391304000000,-0.017211642726301084000000,0.013862497435846789000000,-0.059750627717945648000000,-0.124362460751525470000000,0.197704818771195060000000,0.695739150561516030000000,0.644564383901189420000000,0.110230223021359150000000,-0.140490093113647320000000,0.008819757670415267700000,0.092926030899134981000000,0.017618296880650790000000,-0.020749686325516842000000,-0.001492447274259776600000,0.005674853760122613000000,0.000413261198841939770000,-0.000721364385136249440000,0.000036905373423202441000,0.000070429866906947011000};
localparam real pSYM13_Lo_R [26] = '{0.000070429866906947011000,0.000036905373423202441000,-0.000721364385136249440000,0.000413261198841939770000,0.005674853760122613000000,-0.001492447274259776600000,-0.020749686325516842000000,0.017618296880650790000000,0.092926030899134981000000,0.008819757670415267700000,-0.140490093113647320000000,0.110230223021359150000000,0.644564383901189420000000,0.695739150561516030000000,0.197704818771195060000000,-0.124362460751525470000000,-0.059750627717945648000000,0.013862497435846789000000,-0.017211642726301084000000,-0.020216768133391304000000,0.005296359738724500500000,0.007526225389968108300000,-0.000170942858530178690000,-0.001136063438928119200000,-0.000035738623648692444000,0.000068203252630752971000};
localparam real pSYM13_Hi_D [26] = '{-0.000070429866906947011000,0.000036905373423202441000,0.000721364385136249440000,0.000413261198841939770000,-0.005674853760122613000000,-0.001492447274259776600000,0.020749686325516842000000,0.017618296880650790000000,-0.092926030899134981000000,0.008819757670415267700000,0.140490093113647320000000,0.110230223021359150000000,-0.644564383901189420000000,0.695739150561516030000000,-0.197704818771195060000000,-0.124362460751525470000000,0.059750627717945648000000,0.013862497435846789000000,0.017211642726301084000000,-0.020216768133391304000000,-0.005296359738724500500000,0.007526225389968108300000,0.000170942858530178690000,-0.001136063438928119200000,0.000035738623648692444000,0.000068203252630752971000};
localparam real pSYM13_Hi_R [26] = '{0.000068203252630752971000,0.000035738623648692444000,-0.001136063438928119200000,0.000170942858530178690000,0.007526225389968108300000,-0.005296359738724500500000,-0.020216768133391304000000,0.017211642726301084000000,0.013862497435846789000000,0.059750627717945648000000,-0.124362460751525470000000,-0.197704818771195060000000,0.695739150561516030000000,-0.644564383901189420000000,0.110230223021359150000000,0.140490093113647320000000,0.008819757670415267700000,-0.092926030899134981000000,0.017618296880650790000000,0.020749686325516842000000,-0.001492447274259776600000,-0.005674853760122613000000,0.000413261198841939770000,0.000721364385136249440000,0.000036905373423202441000,-0.000070429866906947011000};

localparam real pSYM14_Lo_D [28] = '{-0.000025879090265409365000,0.000011210865808905823000,0.000398435672976186650000,-0.000062865424814709494000,-0.002579441725934396400000,0.000366476573660040010000,0.010037693717678001000000,-0.002753774791223648700000,-0.029196217764058237000000,0.004280520498995491100000,0.037433088362817647000000,-0.057634498351459444000000,-0.035318112115187240000000,0.393201521962039780000000,0.759976241961305980000000,0.475335762634446100000000,-0.058111823317667580000000,-0.159997411146572070000000,0.025898587531037374000000,0.069827616361827383000000,-0.002365048836737275600000,-0.019439314263632251000000,0.001013141987183896200000,0.004532677471947149500000,-0.000073214213566773824000,-0.000605760182466511090000,0.000019329016965553380000,0.000044618977991492056000};
localparam real pSYM14_Lo_R [28] = '{0.000044618977991492056000,0.000019329016965553380000,-0.000605760182466511090000,-0.000073214213566773824000,0.004532677471947149500000,0.001013141987183896200000,-0.019439314263632251000000,-0.002365048836737275600000,0.069827616361827383000000,0.025898587531037374000000,-0.159997411146572070000000,-0.058111823317667580000000,0.475335762634446100000000,0.759976241961305980000000,0.393201521962039780000000,-0.035318112115187240000000,-0.057634498351459444000000,0.037433088362817647000000,0.004280520498995491100000,-0.029196217764058237000000,-0.002753774791223648700000,0.010037693717678001000000,0.000366476573660040010000,-0.002579441725934396400000,-0.000062865424814709494000,0.000398435672976186650000,0.000011210865808905823000,-0.000025879090265409365000};
localparam real pSYM14_Hi_D [28] = '{-0.000044618977991492056000,0.000019329016965553380000,0.000605760182466511090000,-0.000073214213566773824000,-0.004532677471947149500000,0.001013141987183896200000,0.019439314263632251000000,-0.002365048836737275600000,-0.069827616361827383000000,0.025898587531037374000000,0.159997411146572070000000,-0.058111823317667580000000,-0.475335762634446100000000,0.759976241961305980000000,-0.393201521962039780000000,-0.035318112115187240000000,0.057634498351459444000000,0.037433088362817647000000,-0.004280520498995491100000,-0.029196217764058237000000,0.002753774791223648700000,0.010037693717678001000000,-0.000366476573660040010000,-0.002579441725934396400000,0.000062865424814709494000,0.000398435672976186650000,-0.000011210865808905823000,-0.000025879090265409365000};
localparam real pSYM14_Hi_R [28] = '{-0.000025879090265409365000,-0.000011210865808905823000,0.000398435672976186650000,0.000062865424814709494000,-0.002579441725934396400000,-0.000366476573660040010000,0.010037693717678001000000,0.002753774791223648700000,-0.029196217764058237000000,-0.004280520498995491100000,0.037433088362817647000000,0.057634498351459444000000,-0.035318112115187240000000,-0.393201521962039780000000,0.759976241961305980000000,-0.475335762634446100000000,-0.058111823317667580000000,0.159997411146572070000000,0.025898587531037374000000,-0.069827616361827383000000,-0.002365048836737275600000,0.019439314263632251000000,0.001013141987183896200000,-0.004532677471947149500000,-0.000073214213566773824000,0.000605760182466511090000,0.000019329016965553380000,-0.000044618977991492056000};

localparam real pSYM15_Lo_D [30] = '{0.000009712419737965761900,-0.000007359666798927995800,-0.000160661866375015850000,0.000055122547855632115000,0.001070567219462822800000,-0.000267316446471904940000,-0.003590165447373799200000,0.003423450736352785800000,0.010079977087907843000000,-0.019405011430949529000000,-0.038876716876869652000000,0.021937642719713057000000,0.040735479696734966000000,-0.041082666635527246000000,0.111533695142521830000000,0.578640415215140650000000,0.721843029636393240000000,0.243962705432254210000000,-0.196626358766280760000000,-0.134056298456272540000000,0.068393310060520948000000,0.067969829044907476000000,-0.008744788886480820900000,-0.017171252781644327000000,0.001526138278182918300000,0.003481028737066057700000,-0.000108154401685598040000,-0.000402168537603076480000,0.000021717890150803856000,0.000028660708525331908000};
localparam real pSYM15_Lo_R [30] = '{0.000028660708525331908000,0.000021717890150803856000,-0.000402168537603076480000,-0.000108154401685598040000,0.003481028737066057700000,0.001526138278182918300000,-0.017171252781644327000000,-0.008744788886480820900000,0.067969829044907476000000,0.068393310060520948000000,-0.134056298456272540000000,-0.196626358766280760000000,0.243962705432254210000000,0.721843029636393240000000,0.578640415215140650000000,0.111533695142521830000000,-0.041082666635527246000000,0.040735479696734966000000,0.021937642719713057000000,-0.038876716876869652000000,-0.019405011430949529000000,0.010079977087907843000000,0.003423450736352785800000,-0.003590165447373799200000,-0.000267316446471904940000,0.001070567219462822800000,0.000055122547855632115000,-0.000160661866375015850000,-0.000007359666798927995800,0.000009712419737965761900};
localparam real pSYM15_Hi_D [30] = '{-0.000028660708525331908000,0.000021717890150803856000,0.000402168537603076480000,-0.000108154401685598040000,-0.003481028737066057700000,0.001526138278182918300000,0.017171252781644327000000,-0.008744788886480820900000,-0.067969829044907476000000,0.068393310060520948000000,0.134056298456272540000000,-0.196626358766280760000000,-0.243962705432254210000000,0.721843029636393240000000,-0.578640415215140650000000,0.111533695142521830000000,0.041082666635527246000000,0.040735479696734966000000,-0.021937642719713057000000,-0.038876716876869652000000,0.019405011430949529000000,0.010079977087907843000000,-0.003423450736352785800000,-0.003590165447373799200000,0.000267316446471904940000,0.001070567219462822800000,-0.000055122547855632115000,-0.000160661866375015850000,0.000007359666798927995800,0.000009712419737965761900};
localparam real pSYM15_Hi_R [30] = '{0.000009712419737965761900,0.000007359666798927995800,-0.000160661866375015850000,-0.000055122547855632115000,0.001070567219462822800000,0.000267316446471904940000,-0.003590165447373799200000,-0.003423450736352785800000,0.010079977087907843000000,0.019405011430949529000000,-0.038876716876869652000000,-0.021937642719713057000000,0.040735479696734966000000,0.041082666635527246000000,0.111533695142521830000000,-0.578640415215140650000000,0.721843029636393240000000,-0.243962705432254210000000,-0.196626358766280760000000,0.134056298456272540000000,0.068393310060520948000000,-0.067969829044907476000000,-0.008744788886480820900000,0.017171252781644327000000,0.001526138278182918300000,-0.003481028737066057700000,-0.000108154401685598040000,0.000402168537603076480000,0.000021717890150803856000,-0.000028660708525331908000};

localparam real pSYM16_Lo_D [32] = '{0.000006230006701215267600,-0.000003113556407650880500,-0.000109431479295290120000,0.000028078582128712609000,0.000852354710804932970000,-0.000108445622310089130000,-0.003880912252605258100000,0.000718211978833800540000,0.012666731659854047000000,-0.003126517172303187000000,-0.031051202843619220000000,0.004869274404809647400000,0.032333091610498403000000,-0.066983049070456463000000,-0.034574228417094573000000,0.397122933620832900000000,0.756524987876045050000000,0.475342806011696540000000,-0.054040601387650766000000,-0.159592192185254940000000,0.030721139063339703000000,0.078037852903466848000000,-0.003510275068362536300000,-0.024952758046288760000000,0.001359844742489502200000,0.006937761130805780900000,-0.000222116476211911960000,-0.001338720606692478000000,0.000036565924833582383000,0.000165456795791117920000,-0.000005396483179336830300,-0.000010797982104326530000};
localparam real pSYM16_Lo_R [32] = '{-0.000010797982104326530000,-0.000005396483179336830300,0.000165456795791117920000,0.000036565924833582383000,-0.001338720606692478000000,-0.000222116476211911960000,0.006937761130805780900000,0.001359844742489502200000,-0.024952758046288760000000,-0.003510275068362536300000,0.078037852903466848000000,0.030721139063339703000000,-0.159592192185254940000000,-0.054040601387650766000000,0.475342806011696540000000,0.756524987876045050000000,0.397122933620832900000000,-0.034574228417094573000000,-0.066983049070456463000000,0.032333091610498403000000,0.004869274404809647400000,-0.031051202843619220000000,-0.003126517172303187000000,0.012666731659854047000000,0.000718211978833800540000,-0.003880912252605258100000,-0.000108445622310089130000,0.000852354710804932970000,0.000028078582128712609000,-0.000109431479295290120000,-0.000003113556407650880500,0.000006230006701215267600};
localparam real pSYM16_Hi_D [32] = '{0.000010797982104326530000,-0.000005396483179336830300,-0.000165456795791117920000,0.000036565924833582383000,0.001338720606692478000000,-0.000222116476211911960000,-0.006937761130805780900000,0.001359844742489502200000,0.024952758046288760000000,-0.003510275068362536300000,-0.078037852903466848000000,0.030721139063339703000000,0.159592192185254940000000,-0.054040601387650766000000,-0.475342806011696540000000,0.756524987876045050000000,-0.397122933620832900000000,-0.034574228417094573000000,0.066983049070456463000000,0.032333091610498403000000,-0.004869274404809647400000,-0.031051202843619220000000,0.003126517172303187000000,0.012666731659854047000000,-0.000718211978833800540000,-0.003880912252605258100000,0.000108445622310089130000,0.000852354710804932970000,-0.000028078582128712609000,-0.000109431479295290120000,0.000003113556407650880500,0.000006230006701215267600};
localparam real pSYM16_Hi_R [32] = '{0.000006230006701215267600,0.000003113556407650880500,-0.000109431479295290120000,-0.000028078582128712609000,0.000852354710804932970000,0.000108445622310089130000,-0.003880912252605258100000,-0.000718211978833800540000,0.012666731659854047000000,0.003126517172303187000000,-0.031051202843619220000000,-0.004869274404809647400000,0.032333091610498403000000,0.066983049070456463000000,-0.034574228417094573000000,-0.397122933620832900000000,0.756524987876045050000000,-0.475342806011696540000000,-0.054040601387650766000000,0.159592192185254940000000,0.030721139063339703000000,-0.078037852903466848000000,-0.003510275068362536300000,0.024952758046288760000000,0.001359844742489502200000,-0.006937761130805780900000,-0.000222116476211911960000,0.001338720606692478000000,0.000036565924833582383000,-0.000165456795791117920000,-0.000005396483179336830300,0.000010797982104326530000};

localparam real pSYM17_Lo_D [34] = '{0.000004297343327345718700,0.000002780126693852938500,-0.000062937025975495122000,-0.000013506383399943850000,0.000475996380263645670000,-0.000138642302679820490000,-0.002741675975679997600000,0.000856770070188555130000,0.010482366933024175000000,-0.004819212803168662500000,-0.033291383492347310000000,0.017903952214289105000000,0.104754614842132040000000,0.017271178210522237000000,-0.118566932611364330000000,0.142398350414505270000000,0.650716629204113880000000,0.681488995344720180000000,0.180539584581378140000000,-0.155076005349371940000000,-0.086070874720574411000000,0.016158808725943996000000,-0.007261634750896922200000,-0.018038897241896449000000,0.009952982523502705600000,0.012396988366643208000000,-0.001905407689847316700000,-0.003932325279794507400000,0.000058400428693269492000,0.000719827064214206360000,0.000025207933140917839000,-0.000076071244055967002000,-0.000002452716342590583600,0.000003791253194326478500};
localparam real pSYM17_Lo_R [34] = '{0.000003791253194326478500,-0.000002452716342590583600,-0.000076071244055967002000,0.000025207933140917839000,0.000719827064214206360000,0.000058400428693269492000,-0.003932325279794507400000,-0.001905407689847316700000,0.012396988366643208000000,0.009952982523502705600000,-0.018038897241896449000000,-0.007261634750896922200000,0.016158808725943996000000,-0.086070874720574411000000,-0.155076005349371940000000,0.180539584581378140000000,0.681488995344720180000000,0.650716629204113880000000,0.142398350414505270000000,-0.118566932611364330000000,0.017271178210522237000000,0.104754614842132040000000,0.017903952214289105000000,-0.033291383492347310000000,-0.004819212803168662500000,0.010482366933024175000000,0.000856770070188555130000,-0.002741675975679997600000,-0.000138642302679820490000,0.000475996380263645670000,-0.000013506383399943850000,-0.000062937025975495122000,0.000002780126693852938500,0.000004297343327345718700};
localparam real pSYM17_Hi_D [34] = '{-0.000003791253194326478500,-0.000002452716342590583600,0.000076071244055967002000,0.000025207933140917839000,-0.000719827064214206360000,0.000058400428693269492000,0.003932325279794507400000,-0.001905407689847316700000,-0.012396988366643208000000,0.009952982523502705600000,0.018038897241896449000000,-0.007261634750896922200000,-0.016158808725943996000000,-0.086070874720574411000000,0.155076005349371940000000,0.180539584581378140000000,-0.681488995344720180000000,0.650716629204113880000000,-0.142398350414505270000000,-0.118566932611364330000000,-0.017271178210522237000000,0.104754614842132040000000,-0.017903952214289105000000,-0.033291383492347310000000,0.004819212803168662500000,0.010482366933024175000000,-0.000856770070188555130000,-0.002741675975679997600000,0.000138642302679820490000,0.000475996380263645670000,0.000013506383399943850000,-0.000062937025975495122000,-0.000002780126693852938500,0.000004297343327345718700};
localparam real pSYM17_Hi_R [34] = '{0.000004297343327345718700,-0.000002780126693852938500,-0.000062937025975495122000,0.000013506383399943850000,0.000475996380263645670000,0.000138642302679820490000,-0.002741675975679997600000,-0.000856770070188555130000,0.010482366933024175000000,0.004819212803168662500000,-0.033291383492347310000000,-0.017903952214289105000000,0.104754614842132040000000,-0.017271178210522237000000,-0.118566932611364330000000,-0.142398350414505270000000,0.650716629204113880000000,-0.681488995344720180000000,0.180539584581378140000000,0.155076005349371940000000,-0.086070874720574411000000,-0.016158808725943996000000,-0.007261634750896922200000,0.018038897241896449000000,0.009952982523502705600000,-0.012396988366643208000000,-0.001905407689847316700000,0.003932325279794507400000,0.000058400428693269492000,-0.000719827064214206360000,0.000025207933140917839000,0.000076071244055967002000,-0.000002452716342590583600,-0.000003791253194326478500};

localparam real pSYM18_Lo_D [36] = '{0.000002612612556350492500,0.000001354915761541965200,-0.000045246757873133215000,-0.000014020992573916282000,0.000396168406369346120000,0.000070212734565581930000,-0.002313871814432167000000,-0.000411521109091850440000,0.009502164390753133400000,0.001642986396908572300000,-0.030325091088450135000000,-0.005077085158959507300000,0.084219929969611737000000,0.033995667102118238000000,-0.159938148662873620000000,-0.052029158967992123000000,0.473969059904092600000000,0.753629140095299020000000,0.401483860557063870000000,-0.032480573297721249000000,-0.073799207292583741000000,0.028529597037456399000000,0.006277944553024958000000,-0.031712684731719745000000,-0.003260744199722687500000,0.015012356344109535000000,0.001087784789426010500000,-0.005239789682997976700000,-0.000188776239365721810000,0.001428086327075219400000,0.000047416145174328255000,-0.000265830110241911410000,-0.000009858816029108966500,0.000029557437620941463000,0.000000784729805549380270,-0.000001513153069233471200};
localparam real pSYM18_Lo_R [36] = '{-0.000001513153069233471200,0.000000784729805549380270,0.000029557437620941463000,-0.000009858816029108966500,-0.000265830110241911410000,0.000047416145174328255000,0.001428086327075219400000,-0.000188776239365721810000,-0.005239789682997976700000,0.001087784789426010500000,0.015012356344109535000000,-0.003260744199722687500000,-0.031712684731719745000000,0.006277944553024958000000,0.028529597037456399000000,-0.073799207292583741000000,-0.032480573297721249000000,0.401483860557063870000000,0.753629140095299020000000,0.473969059904092600000000,-0.052029158967992123000000,-0.159938148662873620000000,0.033995667102118238000000,0.084219929969611737000000,-0.005077085158959507300000,-0.030325091088450135000000,0.001642986396908572300000,0.009502164390753133400000,-0.000411521109091850440000,-0.002313871814432167000000,0.000070212734565581930000,0.000396168406369346120000,-0.000014020992573916282000,-0.000045246757873133215000,0.000001354915761541965200,0.000002612612556350492500};
localparam real pSYM18_Hi_D [36] = '{0.000001513153069233471200,0.000000784729805549380270,-0.000029557437620941463000,-0.000009858816029108966500,0.000265830110241911410000,0.000047416145174328255000,-0.001428086327075219400000,-0.000188776239365721810000,0.005239789682997976700000,0.001087784789426010500000,-0.015012356344109535000000,-0.003260744199722687500000,0.031712684731719745000000,0.006277944553024958000000,-0.028529597037456399000000,-0.073799207292583741000000,0.032480573297721249000000,0.401483860557063870000000,-0.753629140095299020000000,0.473969059904092600000000,0.052029158967992123000000,-0.159938148662873620000000,-0.033995667102118238000000,0.084219929969611737000000,0.005077085158959507300000,-0.030325091088450135000000,-0.001642986396908572300000,0.009502164390753133400000,0.000411521109091850440000,-0.002313871814432167000000,-0.000070212734565581930000,0.000396168406369346120000,0.000014020992573916282000,-0.000045246757873133215000,-0.000001354915761541965200,0.000002612612556350492500};
localparam real pSYM18_Hi_R [36] = '{0.000002612612556350492500,-0.000001354915761541965200,-0.000045246757873133215000,0.000014020992573916282000,0.000396168406369346120000,-0.000070212734565581930000,-0.002313871814432167000000,0.000411521109091850440000,0.009502164390753133400000,-0.001642986396908572300000,-0.030325091088450135000000,0.005077085158959507300000,0.084219929969611737000000,-0.033995667102118238000000,-0.159938148662873620000000,0.052029158967992123000000,0.473969059904092600000000,-0.753629140095299020000000,0.401483860557063870000000,0.032480573297721249000000,-0.073799207292583741000000,-0.028529597037456399000000,0.006277944553024958000000,0.031712684731719745000000,-0.003260744199722687500000,-0.015012356344109535000000,0.001087784789426010500000,0.005239789682997976700000,-0.000188776239365721810000,-0.001428086327075219400000,0.000047416145174328255000,0.000265830110241911410000,-0.000009858816029108966500,-0.000029557437620941463000,0.000000784729805549380270,0.000001513153069233471200};

localparam real pSYM19_Lo_D [38] = '{0.000000548773276806204780,-0.000000646365130355436200,-0.000011880518269510527000,0.000008873312174298990500,0.000115539233333357400000,-0.000046120396007574042000,-0.000635764514995112560000,0.000159158047705974330000,0.002121425028165130500000,-0.001160703257238153000000,-0.005122205002453399800000,0.007968438320719886000000,0.015797439295212053000000,-0.022651993378824325000000,-0.046635983534439242000000,0.007015573858210684600000,0.008954591174112291900000,-0.067525058035497368000000,0.109025825091803070000000,0.578144945346146240000000,0.719555525710884660000000,0.258266169223859640000000,-0.176596866259597890000000,-0.116241730106131410000000,0.093630843418263096000000,0.084072676278559993000000,-0.016908234862673219000000,-0.027709896931392881000000,0.004319351875256709000000,0.008262236955576022000000,-0.000617922327885841330000,-0.001704960261181416900000,0.000129307676522794170000,0.000276218776860900430000,-0.000016821387031260756000,-0.000028151138661953039000,0.000002062317063419342600,0.000001750936799581956800};
localparam real pSYM19_Lo_R [38] = '{0.000001750936799581956800,0.000002062317063419342600,-0.000028151138661953039000,-0.000016821387031260756000,0.000276218776860900430000,0.000129307676522794170000,-0.001704960261181416900000,-0.000617922327885841330000,0.008262236955576022000000,0.004319351875256709000000,-0.027709896931392881000000,-0.016908234862673219000000,0.084072676278559993000000,0.093630843418263096000000,-0.116241730106131410000000,-0.176596866259597890000000,0.258266169223859640000000,0.719555525710884660000000,0.578144945346146240000000,0.109025825091803070000000,-0.067525058035497368000000,0.008954591174112291900000,0.007015573858210684600000,-0.046635983534439242000000,-0.022651993378824325000000,0.015797439295212053000000,0.007968438320719886000000,-0.005122205002453399800000,-0.001160703257238153000000,0.002121425028165130500000,0.000159158047705974330000,-0.000635764514995112560000,-0.000046120396007574042000,0.000115539233333357400000,0.000008873312174298990500,-0.000011880518269510527000,-0.000000646365130355436200,0.000000548773276806204780};
localparam real pSYM19_Hi_D [38] = '{-0.000001750936799581956800,0.000002062317063419342600,0.000028151138661953039000,-0.000016821387031260756000,-0.000276218776860900430000,0.000129307676522794170000,0.001704960261181416900000,-0.000617922327885841330000,-0.008262236955576022000000,0.004319351875256709000000,0.027709896931392881000000,-0.016908234862673219000000,-0.084072676278559993000000,0.093630843418263096000000,0.116241730106131410000000,-0.176596866259597890000000,-0.258266169223859640000000,0.719555525710884660000000,-0.578144945346146240000000,0.109025825091803070000000,0.067525058035497368000000,0.008954591174112291900000,-0.007015573858210684600000,-0.046635983534439242000000,0.022651993378824325000000,0.015797439295212053000000,-0.007968438320719886000000,-0.005122205002453399800000,0.001160703257238153000000,0.002121425028165130500000,-0.000159158047705974330000,-0.000635764514995112560000,0.000046120396007574042000,0.000115539233333357400000,-0.000008873312174298990500,-0.000011880518269510527000,0.000000646365130355436200,0.000000548773276806204780};
localparam real pSYM19_Hi_R [38] = '{0.000000548773276806204780,0.000000646365130355436200,-0.000011880518269510527000,-0.000008873312174298990500,0.000115539233333357400000,0.000046120396007574042000,-0.000635764514995112560000,-0.000159158047705974330000,0.002121425028165130500000,0.001160703257238153000000,-0.005122205002453399800000,-0.007968438320719886000000,0.015797439295212053000000,0.022651993378824325000000,-0.046635983534439242000000,-0.007015573858210684600000,0.008954591174112291900000,0.067525058035497368000000,0.109025825091803070000000,-0.578144945346146240000000,0.719555525710884660000000,-0.258266169223859640000000,-0.176596866259597890000000,0.116241730106131410000000,0.093630843418263096000000,-0.084072676278559993000000,-0.016908234862673219000000,0.027709896931392881000000,0.004319351875256709000000,-0.008262236955576022000000,-0.000617922327885841330000,0.001704960261181416900000,0.000129307676522794170000,-0.000276218776860900430000,-0.000016821387031260756000,0.000028151138661953039000,0.000002062317063419342600,-0.000001750936799581956800};

localparam real pSYM20_Lo_D [40] = '{0.000000369553747499528320,-0.000000190156758914925810,-0.000007919361412311997100,0.000003025666062914772300,0.000079929678361088981000,-0.000019284123007819317000,-0.000494731091588121730000,0.000072159911886191406000,0.002088994708271114300000,-0.000305262831846022230000,-0.006606585799414299400000,0.001423087359477369700000,0.017004049023916480000000,-0.003313857384204183600000,-0.031629437146754244000000,0.008123228355724163400000,0.025579349508645426000000,-0.078994344935197788000000,-0.029819368885983914000000,0.405831444358891070000000,0.751162728442403950000000,0.471991475106061820000000,-0.051088342934149843000000,-0.160578298424811470000000,0.036250951656373251000000,0.088919668031744795000000,-0.006843701966416111000000,-0.035373336758335407000000,0.001938597067621526000000,0.012157040949352209000000,-0.000611126385943504400000,-0.003471647803017408700000,0.000125440917266307330000,0.000747610859821253700000,-0.000026615550342593026000,-0.000117391335169443810000,0.000004525422210144222400,0.000012287252778689056000,-0.000000325670264284955790,-0.000000632912904524793580};
localparam real pSYM20_Lo_R [40] = '{-0.000000632912904524793580,-0.000000325670264284955790,0.000012287252778689056000,0.000004525422210144222400,-0.000117391335169443810000,-0.000026615550342593026000,0.000747610859821253700000,0.000125440917266307330000,-0.003471647803017408700000,-0.000611126385943504400000,0.012157040949352209000000,0.001938597067621526000000,-0.035373336758335407000000,-0.006843701966416111000000,0.088919668031744795000000,0.036250951656373251000000,-0.160578298424811470000000,-0.051088342934149843000000,0.471991475106061820000000,0.751162728442403950000000,0.405831444358891070000000,-0.029819368885983914000000,-0.078994344935197788000000,0.025579349508645426000000,0.008123228355724163400000,-0.031629437146754244000000,-0.003313857384204183600000,0.017004049023916480000000,0.001423087359477369700000,-0.006606585799414299400000,-0.000305262831846022230000,0.002088994708271114300000,0.000072159911886191406000,-0.000494731091588121730000,-0.000019284123007819317000,0.000079929678361088981000,0.000003025666062914772300,-0.000007919361412311997100,-0.000000190156758914925810,0.000000369553747499528320};
localparam real pSYM20_Hi_D [40] = '{0.000000632912904524793580,-0.000000325670264284955790,-0.000012287252778689056000,0.000004525422210144222400,0.000117391335169443810000,-0.000026615550342593026000,-0.000747610859821253700000,0.000125440917266307330000,0.003471647803017408700000,-0.000611126385943504400000,-0.012157040949352209000000,0.001938597067621526000000,0.035373336758335407000000,-0.006843701966416111000000,-0.088919668031744795000000,0.036250951656373251000000,0.160578298424811470000000,-0.051088342934149843000000,-0.471991475106061820000000,0.751162728442403950000000,-0.405831444358891070000000,-0.029819368885983914000000,0.078994344935197788000000,0.025579349508645426000000,-0.008123228355724163400000,-0.031629437146754244000000,0.003313857384204183600000,0.017004049023916480000000,-0.001423087359477369700000,-0.006606585799414299400000,0.000305262831846022230000,0.002088994708271114300000,-0.000072159911886191406000,-0.000494731091588121730000,0.000019284123007819317000,0.000079929678361088981000,-0.000003025666062914772300,-0.000007919361412311997100,0.000000190156758914925810,0.000000369553747499528320};
localparam real pSYM20_Hi_R [40] = '{0.000000369553747499528320,0.000000190156758914925810,-0.000007919361412311997100,-0.000003025666062914772300,0.000079929678361088981000,0.000019284123007819317000,-0.000494731091588121730000,-0.000072159911886191406000,0.002088994708271114300000,0.000305262831846022230000,-0.006606585799414299400000,-0.001423087359477369700000,0.017004049023916480000000,0.003313857384204183600000,-0.031629437146754244000000,-0.008123228355724163400000,0.025579349508645426000000,0.078994344935197788000000,-0.029819368885983914000000,-0.405831444358891070000000,0.751162728442403950000000,-0.471991475106061820000000,-0.051088342934149843000000,0.160578298424811470000000,0.036250951656373251000000,-0.088919668031744795000000,-0.006843701966416111000000,0.035373336758335407000000,0.001938597067621526000000,-0.012157040949352209000000,-0.000611126385943504400000,0.003471647803017408700000,0.000125440917266307330000,-0.000747610859821253700000,-0.000026615550342593026000,0.000117391335169443810000,0.000004525422210144222400,-0.000012287252778689056000,-0.000000325670264284955790,0.000000632912904524793580};

localparam real pDMEY_Lo_D [102] = '{0.000000000000000000000000,-0.000001509740857423615400,0.000001278766756823498800,0.000000449585560448868940,-0.000002096568870494942400,0.000001723223554480681600,0.000000698082276310738600,-0.000002879408032654846900,0.000002383148394518929800,0.000000982515602229338580,-0.000004217789186342479200,0.000003353501538089443700,0.000001674721858836507200,-0.000006034501341860346700,0.000004837555801559578900,0.000002402288022882837700,-0.000009556309845665444700,0.000007216527694763414900,0.000004849078299776748700,-0.000014206928580564191000,0.000010503914270783866000,0.000006187580298111554400,-0.000024438005845654610000,0.000020106387690909483000,0.000014993523600015134000,-0.000046428764283651690000,0.000032341311913679687000,0.000037409665760249841000,-0.000102779005084884770000,0.000024461956844602302000,0.000149713515389257360000,-0.000075592870255167127000,-0.000139913148217418020000,-0.000093512893880113803000,0.000161189819725346310000,0.000859500213762377500000,-0.000578185795273441120000,-0.002702168733939079700000,0.002194775336459444400000,0.006045510596456077700000,-0.006386728618548126300000,-0.011044641900538889000000,0.015250913158585904000000,0.017403888210177406000000,-0.032094063354505306000000,-0.024321783959518777000000,0.063667300884468314000000,0.030621243943424570000000,-0.132696615358861740000000,-0.035048287390595033000000,0.444095030766528790000000,0.743751004903786980000000,0.444095030766528790000000,-0.035048287390595033000000,-0.132696615358861740000000,0.030621243943424570000000,0.063667300884468314000000,-0.024321783959518777000000,-0.032094063354505306000000,0.017403888210177406000000,0.015250913158585904000000,-0.011044641900538889000000,-0.006386728618548126300000,0.006045510596456077700000,0.002194775336459444400000,-0.002702168733939079700000,-0.000578185795273441120000,0.000859500213762377500000,0.000161189819725346310000,-0.000093512893880113803000,-0.000139913148217418020000,-0.000075592870255167127000,0.000149713515389257360000,0.000024461956844602302000,-0.000102779005084884770000,0.000037409665760249841000,0.000032341311913679687000,-0.000046428764283651690000,0.000014993523600015134000,0.000020106387690909483000,-0.000024438005845654610000,0.000006187580298111554400,0.000010503914270783866000,-0.000014206928580564191000,0.000004849078299776748700,0.000007216527694763414900,-0.000009556309845665444700,0.000002402288022882837700,0.000004837555801559578900,-0.000006034501341860346700,0.000001674721858836507200,0.000003353501538089443700,-0.000004217789186342479200,0.000000982515602229338580,0.000002383148394518929800,-0.000002879408032654846900,0.000000698082276310738600,0.000001723223554480681600,-0.000002096568870494942400,0.000000449585560448868940,0.000001278766756823498800,-0.000001509740857423615400};
localparam real pDMEY_Lo_R [102] = '{-0.000001509740857423615400,0.000001278766756823498800,0.000000449585560448868940,-0.000002096568870494942400,0.000001723223554480681600,0.000000698082276310738600,-0.000002879408032654846900,0.000002383148394518929800,0.000000982515602229338580,-0.000004217789186342479200,0.000003353501538089443700,0.000001674721858836507200,-0.000006034501341860346700,0.000004837555801559578900,0.000002402288022882837700,-0.000009556309845665444700,0.000007216527694763414900,0.000004849078299776748700,-0.000014206928580564191000,0.000010503914270783866000,0.000006187580298111554400,-0.000024438005845654610000,0.000020106387690909483000,0.000014993523600015134000,-0.000046428764283651690000,0.000032341311913679687000,0.000037409665760249841000,-0.000102779005084884770000,0.000024461956844602302000,0.000149713515389257360000,-0.000075592870255167127000,-0.000139913148217418020000,-0.000093512893880113803000,0.000161189819725346310000,0.000859500213762377500000,-0.000578185795273441120000,-0.002702168733939079700000,0.002194775336459444400000,0.006045510596456077700000,-0.006386728618548126300000,-0.011044641900538889000000,0.015250913158585904000000,0.017403888210177406000000,-0.032094063354505306000000,-0.024321783959518777000000,0.063667300884468314000000,0.030621243943424570000000,-0.132696615358861740000000,-0.035048287390595033000000,0.444095030766528790000000,0.743751004903786980000000,0.444095030766528790000000,-0.035048287390595033000000,-0.132696615358861740000000,0.030621243943424570000000,0.063667300884468314000000,-0.024321783959518777000000,-0.032094063354505306000000,0.017403888210177406000000,0.015250913158585904000000,-0.011044641900538889000000,-0.006386728618548126300000,0.006045510596456077700000,0.002194775336459444400000,-0.002702168733939079700000,-0.000578185795273441120000,0.000859500213762377500000,0.000161189819725346310000,-0.000093512893880113803000,-0.000139913148217418020000,-0.000075592870255167127000,0.000149713515389257360000,0.000024461956844602302000,-0.000102779005084884770000,0.000037409665760249841000,0.000032341311913679687000,-0.000046428764283651690000,0.000014993523600015134000,0.000020106387690909483000,-0.000024438005845654610000,0.000006187580298111554400,0.000010503914270783866000,-0.000014206928580564191000,0.000004849078299776748700,0.000007216527694763414900,-0.000009556309845665444700,0.000002402288022882837700,0.000004837555801559578900,-0.000006034501341860346700,0.000001674721858836507200,0.000003353501538089443700,-0.000004217789186342479200,0.000000982515602229338580,0.000002383148394518929800,-0.000002879408032654846900,0.000000698082276310738600,0.000001723223554480681600,-0.000002096568870494942400,0.000000449585560448868940,0.000001278766756823498800,-0.000001509740857423615400,0.000000000000000000000000};
localparam real pDMEY_Hi_D [102] = '{0.000001509740857423615400,0.000001278766756823498800,-0.000000449585560448868940,-0.000002096568870494942400,-0.000001723223554480681600,0.000000698082276310738600,0.000002879408032654846900,0.000002383148394518929800,-0.000000982515602229338580,-0.000004217789186342479200,-0.000003353501538089443700,0.000001674721858836507200,0.000006034501341860346700,0.000004837555801559578900,-0.000002402288022882837700,-0.000009556309845665444700,-0.000007216527694763414900,0.000004849078299776748700,0.000014206928580564191000,0.000010503914270783866000,-0.000006187580298111554400,-0.000024438005845654610000,-0.000020106387690909483000,0.000014993523600015134000,0.000046428764283651690000,0.000032341311913679687000,-0.000037409665760249841000,-0.000102779005084884770000,-0.000024461956844602302000,0.000149713515389257360000,0.000075592870255167127000,-0.000139913148217418020000,0.000093512893880113803000,0.000161189819725346310000,-0.000859500213762377500000,-0.000578185795273441120000,0.002702168733939079700000,0.002194775336459444400000,-0.006045510596456077700000,-0.006386728618548126300000,0.011044641900538889000000,0.015250913158585904000000,-0.017403888210177406000000,-0.032094063354505306000000,0.024321783959518777000000,0.063667300884468314000000,-0.030621243943424570000000,-0.132696615358861740000000,0.035048287390595033000000,0.444095030766528790000000,-0.743751004903786980000000,0.444095030766528790000000,0.035048287390595033000000,-0.132696615358861740000000,-0.030621243943424570000000,0.063667300884468314000000,0.024321783959518777000000,-0.032094063354505306000000,-0.017403888210177406000000,0.015250913158585904000000,0.011044641900538889000000,-0.006386728618548126300000,-0.006045510596456077700000,0.002194775336459444400000,0.002702168733939079700000,-0.000578185795273441120000,-0.000859500213762377500000,0.000161189819725346310000,0.000093512893880113803000,-0.000139913148217418020000,0.000075592870255167127000,0.000149713515389257360000,-0.000024461956844602302000,-0.000102779005084884770000,-0.000037409665760249841000,0.000032341311913679687000,0.000046428764283651690000,0.000014993523600015134000,-0.000020106387690909483000,-0.000024438005845654610000,-0.000006187580298111554400,0.000010503914270783866000,0.000014206928580564191000,0.000004849078299776748700,-0.000007216527694763414900,-0.000009556309845665444700,-0.000002402288022882837700,0.000004837555801559578900,0.000006034501341860346700,0.000001674721858836507200,-0.000003353501538089443700,-0.000004217789186342479200,-0.000000982515602229338580,0.000002383148394518929800,0.000002879408032654846900,0.000000698082276310738600,-0.000001723223554480681600,-0.000002096568870494942400,-0.000000449585560448868940,0.000001278766756823498800,0.000001509740857423615400,0.000000000000000000000000};
localparam real pDMEY_Hi_R [102] = '{0.000000000000000000000000,0.000001509740857423615400,0.000001278766756823498800,-0.000000449585560448868940,-0.000002096568870494942400,-0.000001723223554480681600,0.000000698082276310738600,0.000002879408032654846900,0.000002383148394518929800,-0.000000982515602229338580,-0.000004217789186342479200,-0.000003353501538089443700,0.000001674721858836507200,0.000006034501341860346700,0.000004837555801559578900,-0.000002402288022882837700,-0.000009556309845665444700,-0.000007216527694763414900,0.000004849078299776748700,0.000014206928580564191000,0.000010503914270783866000,-0.000006187580298111554400,-0.000024438005845654610000,-0.000020106387690909483000,0.000014993523600015134000,0.000046428764283651690000,0.000032341311913679687000,-0.000037409665760249841000,-0.000102779005084884770000,-0.000024461956844602302000,0.000149713515389257360000,0.000075592870255167127000,-0.000139913148217418020000,0.000093512893880113803000,0.000161189819725346310000,-0.000859500213762377500000,-0.000578185795273441120000,0.002702168733939079700000,0.002194775336459444400000,-0.006045510596456077700000,-0.006386728618548126300000,0.011044641900538889000000,0.015250913158585904000000,-0.017403888210177406000000,-0.032094063354505306000000,0.024321783959518777000000,0.063667300884468314000000,-0.030621243943424570000000,-0.132696615358861740000000,0.035048287390595033000000,0.444095030766528790000000,-0.743751004903786980000000,0.444095030766528790000000,0.035048287390595033000000,-0.132696615358861740000000,-0.030621243943424570000000,0.063667300884468314000000,0.024321783959518777000000,-0.032094063354505306000000,-0.017403888210177406000000,0.015250913158585904000000,0.011044641900538889000000,-0.006386728618548126300000,-0.006045510596456077700000,0.002194775336459444400000,0.002702168733939079700000,-0.000578185795273441120000,-0.000859500213762377500000,0.000161189819725346310000,0.000093512893880113803000,-0.000139913148217418020000,0.000075592870255167127000,0.000149713515389257360000,-0.000024461956844602302000,-0.000102779005084884770000,-0.000037409665760249841000,0.000032341311913679687000,0.000046428764283651690000,0.000014993523600015134000,-0.000020106387690909483000,-0.000024438005845654610000,-0.000006187580298111554400,0.000010503914270783866000,0.000014206928580564191000,0.000004849078299776748700,-0.000007216527694763414900,-0.000009556309845665444700,-0.000002402288022882837700,0.000004837555801559578900,0.000006034501341860346700,0.000001674721858836507200,-0.000003353501538089443700,-0.000004217789186342479200,-0.000000982515602229338580,0.000002383148394518929800,0.000002879408032654846900,0.000000698082276310738600,-0.000001723223554480681600,-0.000002096568870494942400,-0.000000449585560448868940,0.000001278766756823498800,0.000001509740857423615400};

`endif
