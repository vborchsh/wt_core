
`ifndef __WT_HEADER__
`define __WT_HEADER__

//--------------------------------------------------------------------------------------------------------
// File connection
//--------------------------------------------------------------------------------------------------------

`include "./header_wavelets.svh"
//
`include "./../rtl/wt_common/wt_fir.sv"

//--------------------------------------------------------------------------------------------------------
// Parameters
//--------------------------------------------------------------------------------------------------------

localparam int pW_C                    = 8;
localparam int pC_MULT                 = 2**8;

`endif

