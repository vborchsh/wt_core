localparam bit [15:0] pHAAR_Lo_D [2] = '{23170,23170};
localparam bit [15:0] pHAAR_Lo_R [2] = '{23170,23170};
localparam bit [15:0] pHAAR_Hi_D [2] = '{-23171,23170};
localparam bit [15:0] pHAAR_Hi_R [2] = '{23170,-23171};

localparam bit [15:0] pDB1_Lo_D [2] = '{23170,23170};
localparam bit [15:0] pDB1_Lo_R [2] = '{23170,23170};
localparam bit [15:0] pDB1_Hi_D [2] = '{-23171,23170};
localparam bit [15:0] pDB1_Hi_R [2] = '{23170,-23171};

localparam bit [15:0] pDB2_Lo_D [4] = '{-4241,7344,27410,15825};
localparam bit [15:0] pDB2_Lo_R [4] = '{15825,27410,7344,-4241};
localparam bit [15:0] pDB2_Hi_D [4] = '{-15826,27410,-7345,-4241};
localparam bit [15:0] pDB2_Hi_R [4] = '{-4241,-7345,27410,-15826};

localparam bit [15:0] pDB3_Lo_D [6] = '{1154,-2800,-4425,15069,26440,10900};
localparam bit [15:0] pDB3_Lo_R [6] = '{10900,26440,15069,-4425,-2800,1154};
localparam bit [15:0] pDB3_Hi_D [6] = '{-10901,26440,-15070,-4425,2799,1154};
localparam bit [15:0] pDB3_Hi_R [6] = '{1154,2799,-4425,-15070,26440,-10901};

localparam bit [15:0] pDB4_Lo_D [8] = '{-348,1077,1010,-6129,-917,20672,23424,7549};
localparam bit [15:0] pDB4_Lo_R [8] = '{7549,23424,20672,-917,-6129,1010,1077,-348};
localparam bit [15:0] pDB4_Hi_D [8] = '{-7550,23424,-20673,-917,6128,1010,-1078,-348};
localparam bit [15:0] pDB4_Hi_R [8] = '{-348,-1078,1010,6128,-917,-20673,23424,-7550};

localparam bit [15:0] pDB5_Lo_D [10] = '{109,-413,-205,2541,-1057,-7940,4536,23734,19786,5246};
localparam bit [15:0] pDB5_Lo_R [10] = '{5246,19786,23734,4536,-7940,-1057,2541,-205,-413,109};
localparam bit [15:0] pDB5_Hi_D [10] = '{-5247,19786,-23735,4536,7939,-1057,-2542,-205,412,109};
localparam bit [15:0] pDB5_Hi_R [10] = '{109,412,-205,-2542,-1057,7939,4536,-23735,19786,-5247};

localparam bit [15:0] pDB6_Lo_D [12] = '{-36,156,18,-1035,901,3194,-4253,-7415,10330,24613,16207,3654};
localparam bit [15:0] pDB6_Lo_R [12] = '{3654,16207,24613,10330,-7415,-4253,3194,901,-1035,18,156,-36};
localparam bit [15:0] pDB6_Hi_D [12] = '{-3655,16207,-24614,10330,7414,-4253,-3195,901,1034,18,-157,-36};
localparam bit [15:0] pDB6_Hi_R [12] = '{-36,-157,18,1034,901,-3195,-4253,7414,10330,-24614,16207,-3655};

localparam bit [15:0] pDB7_Lo_D [14] = '{11,-60,14,411,-544,-1247,2641,2336,-7342,-4716,15393,23892,12993,2551};
localparam bit [15:0] pDB7_Lo_R [14] = '{2551,12993,23892,15393,-4716,-7342,2336,2641,-1247,-544,411,14,-60,11};
localparam bit [15:0] pDB7_Hi_D [14] = '{-2552,12993,-23893,15393,4715,-7342,-2337,2641,1246,-544,-412,14,59,11};
localparam bit [15:0] pDB7_Hi_R [14] = '{11,59,14,-412,-544,1246,2641,-2337,-7342,4715,15393,-23893,12993,-2552};

localparam bit [15:0] pDB8_Lo_D [16] = '{-4,22,-13,-160,286,458,-1445,-570,4218,15,-9307,-519,19180,22139,10252,1783};
localparam bit [15:0] pDB8_Lo_R [16] = '{1783,10252,22139,19180,-519,-9307,15,4218,-570,-1445,458,286,-160,-13,22,-4};
localparam bit [15:0] pDB8_Hi_D [16] = '{-1784,10252,-22140,19180,518,-9307,-16,4218,569,-1445,-459,286,159,-13,-23,-4};
localparam bit [15:0] pDB8_Hi_R [16] = '{-4,-23,-13,159,286,-459,-1445,569,4218,-16,-9307,518,19180,-22140,10252,-1784};

localparam bit [15:0] pDB9_Lo_D [18] = '{1,-9,7,60,-141,-155,732,8,-2217,1006,4867,-3174,-9610,4364,21538,19818,7989,1247};
localparam bit [15:0] pDB9_Lo_R [18] = '{1247,7989,19818,21538,4364,-9610,-3174,4867,1006,-2217,8,732,-155,-141,60,7,-9,1};
localparam bit [15:0] pDB9_Hi_D [18] = '{-1248,7989,-19819,21538,-4365,-9610,3173,4867,-1007,-2217,-9,732,154,-141,-61,7,8,1};
localparam bit [15:0] pDB9_Hi_R [18] = '{1,8,7,-61,-141,154,732,-9,-2217,-1007,4867,3173,-9610,-4365,21538,-19819,7989,-1248};

localparam bit [15:0] pDB10_Lo_D [20] = '{-1,3,-4,-23,65,45,-352,118,1088,-966,-2340,3049,4173,-6421,-8187,9213,22559,17275,6166,873};
localparam bit [15:0] pDB10_Lo_R [20] = '{873,6166,17275,22559,9213,-8187,-6421,4173,3049,-2340,-966,1088,118,-352,45,65,-23,-4,3,-1};
localparam bit [15:0] pDB10_Hi_D [20] = '{-874,6166,-17276,22559,-9214,-8187,6420,4173,-3050,-2340,965,1088,-119,-352,-46,65,22,-4,-4,-1};
localparam bit [15:0] pDB10_Hi_R [20] = '{-1,-4,-4,22,65,-46,-352,-119,1088,965,-2340,-3050,4173,6420,-8187,-9214,22559,-17276,6166,-874};

localparam bit [15:0] pDB11_Lo_D [22] = '{0,-2,1,8,-30,-11,161,-110,-504,682,1026,-2178,-1524,4909,2164,-8986,-5318,13499,22468,14742,4720,612};
localparam bit [15:0] pDB11_Lo_R [22] = '{612,4720,14742,22468,13499,-5318,-8986,2164,4909,-1524,-2178,1026,682,-504,-110,161,-11,-30,8,1,-2,0};
localparam bit [15:0] pDB11_Hi_D [22] = '{-613,4720,-14743,22468,-13500,-5318,8985,2164,-4910,-1524,2177,1026,-683,-504,109,161,10,-30,-9,1,1,0};
localparam bit [15:0] pDB11_Hi_R [22] = '{0,1,1,-9,-30,10,161,109,-504,-683,1026,2177,-1524,-4910,2164,8985,-5318,-13500,22468,-14743,4720,-613};

localparam bit [15:0] pDB12_Lo_D [24] = '{-1,0,-1,-3,12,0,-72,73,219,-421,-401,1361,355,-3160,175,5979,-780,-10361,-1467,16904,21535,12365,3590,429};
localparam bit [15:0] pDB12_Lo_R [24] = '{429,3590,12365,21535,16904,-1467,-10361,-780,5979,175,-3160,355,1361,-401,-421,219,73,-72,0,12,-3,-1,0,-1};
localparam bit [15:0] pDB12_Hi_D [24] = '{-430,3590,-12366,21535,-16905,-1467,10360,-780,-5980,175,3159,355,-1362,-401,420,219,-74,-72,-1,12,2,-1,-1,-1};
localparam bit [15:0] pDB12_Hi_R [24] = '{-1,-1,-1,2,12,-1,-72,-74,219,420,-401,-1362,355,3159,175,-5980,-780,10360,-1467,-16905,21535,-12366,3590,-430};

localparam bit [15:0] pDB13_Lo_D [26] = '{0,-1,0,1,-6,1,30,-44,-91,237,128,-781,77,1839,-868,-3468,2390,5881,-4083,-10322,2850,19296,20023,10223,2715,301};
localparam bit [15:0] pDB13_Lo_R [26] = '{301,2715,10223,20023,19296,2850,-10322,-4083,5881,2390,-3468,-868,1839,77,-781,128,237,-91,-44,30,1,-6,1,0,-1,0};
localparam bit [15:0] pDB13_Hi_D [26] = '{-302,2715,-10224,20023,-19297,2850,10321,-4083,-5882,2390,3467,-868,-1840,77,780,128,-238,-91,43,30,-2,-6,-2,0,0,0};
localparam bit [15:0] pDB13_Hi_R [26] = '{0,0,0,-2,-6,-2,30,43,-91,-238,128,780,77,-1840,-868,3467,2390,-5882,-4083,10321,2850,-19297,20023,-10224,2715,-302};

localparam bit [15:0] pDB14_Lo_D [28] = '{-1,0,-1,-1,2,-2,-13,23,34,-127,-25,419,-184,-990,884,1810,-2345,-2843,4587,4534,-7145,-8903,7165,20682,18163,8350,2043,211};
localparam bit [15:0] pDB14_Lo_R [28] = '{211,2043,8350,18163,20682,7165,-8903,-7145,4534,4587,-2843,-2345,1810,884,-990,-184,419,-25,-127,34,23,-13,-2,2,-1,-1,0,-1};
localparam bit [15:0] pDB14_Hi_D [28] = '{-212,2043,-8351,18163,-20683,7165,8902,-7145,-4535,4587,2842,-2345,-1811,884,989,-184,-420,-25,126,34,-24,-13,1,2,0,-1,-1,-1};
localparam bit [15:0] pDB14_Hi_R [28] = '{-1,-1,-1,0,2,1,-13,-24,34,126,-25,-420,-184,989,884,-1811,-2345,2842,4587,-4535,-7145,8902,7165,-20683,18163,-8351,2043,-212};

localparam bit [15:0] pDB15_Lo_D [30] = '{0,-1,0,0,-1,0,5,-12,-13,63,-8,-213,167,494,-682,-845,1795,1110,-3642,-1300,6230,2139,-9467,-6331,11108,21162,16142,6750,1531,148};
localparam bit [15:0] pDB15_Lo_R [30] = '{148,1531,6750,16142,21162,11108,-6331,-9467,2139,6230,-1300,-3642,1110,1795,-845,-682,494,167,-213,-8,63,-13,-12,5,0,-1,0,0,-1,0};
localparam bit [15:0] pDB15_Hi_D [30] = '{-149,1531,-6751,16142,-21163,11108,6330,-9467,-2140,6230,1299,-3642,-1111,1795,844,-682,-495,167,212,-8,-64,-13,11,5,-1,-1,-1,0,0,0};
localparam bit [15:0] pDB15_Hi_R [30] = '{0,0,0,-1,-1,-1,5,11,-13,-64,-8,212,167,-495,-682,844,1795,-1111,-3642,1299,6230,-2140,-9467,6330,11108,-21163,16142,-6751,1531,-149};

localparam bit [15:0] pDB16_Lo_D [32] = '{-1,0,-1,-1,0,-1,-3,5,3,-31,13,102,-120,-230,458,337,-1209,-249,2487,-205,-4339,895,6920,-915,-10718,-2941,14427,20884,14100,5408,1143,104};
localparam bit [15:0] pDB16_Lo_R [32] = '{104,1143,5408,14100,20884,14427,-2941,-10718,-915,6920,895,-4339,-205,2487,-249,-1209,337,458,-230,-120,102,13,-31,3,5,-3,-1,0,-1,-1,0,-1};
localparam bit [15:0] pDB16_Hi_D [32] = '{-105,1143,-5409,14100,-20885,14427,2940,-10718,914,6920,-896,-4339,204,2487,248,-1209,-338,458,229,-120,-103,13,30,3,-6,-3,0,0,0,-1,-1,-1};
localparam bit [15:0] pDB16_Hi_R [32] = '{-1,-1,-1,0,0,0,-3,-6,3,30,13,-103,-120,229,458,-338,-1209,248,2487,204,-4339,-896,6920,914,-10718,2940,14427,-20885,14100,-5409,1143,-105};

localparam bit [15:0] pDB17_Lo_D [34] = '{0,-1,0,0,-1,0,0,-3,-1,14,-11,-48,75,97,-282,-100,744,-108,-1538,731,2657,-1871,-4156,3314,6465,-4149,-10759,895,16984,20021,12135,4299,851,73};
localparam bit [15:0] pDB17_Lo_R [34] = '{73,851,4299,12135,20021,16984,895,-10759,-4149,6465,3314,-4156,-1871,2657,731,-1538,-108,744,-100,-282,97,75,-48,-11,14,-1,-3,0,0,-1,0,0,-1,0};
localparam bit [15:0] pDB17_Hi_D [34] = '{-74,851,-4300,12135,-20022,16984,-896,-10759,4148,6465,-3315,-4156,1870,2657,-732,-1538,107,744,99,-282,-98,75,47,-11,-15,-1,2,0,-1,-1,-1,0,0,0};
localparam bit [15:0] pDB17_Hi_R [34] = '{0,0,0,-1,-1,-1,0,2,-1,-15,-11,47,75,-98,-282,99,744,107,-1538,-732,2657,1870,-4156,-3315,6465,4148,-10759,-896,16984,-20022,12135,-4300,851,-74};

localparam bit [15:0] pDB18_Lo_D [36] = '{-1,0,-1,-1,0,-1,-1,1,-1,-7,6,20,-44,-37,161,3,-428,205,873,-778,-1460,1869,2126,-3499,-3026,5474,4899,-7094,-9623,4824,18736,18737,10311,3394,632,51};
localparam bit [15:0] pDB18_Lo_R [36] = '{51,632,3394,10311,18737,18736,4824,-9623,-7094,4899,5474,-3026,-3499,2126,1869,-1460,-778,873,205,-428,3,161,-37,-44,20,6,-7,-1,1,-1,-1,0,-1,-1,0,-1};
localparam bit [15:0] pDB18_Hi_D [36] = '{-52,632,-3395,10311,-18738,18736,-4825,-9623,7093,4899,-5475,-3026,3498,2126,-1870,-1460,777,873,-206,-428,-4,161,36,-44,-21,6,6,-1,-2,-1,0,0,0,-1,-1,-1};
localparam bit [15:0] pDB18_Hi_R [36] = '{-1,-1,-1,0,0,0,-1,-2,-1,6,6,-21,-44,36,161,-4,-428,-206,873,777,-1460,-1870,2126,3498,-3026,-5475,4899,7093,-9623,-4825,18736,-18738,10311,-3395,632,-52};

localparam bit [15:0] pDB19_Lo_D [38] = '{0,-1,0,0,-1,0,0,-1,0,2,-5,-9,24,11,-89,25,230,-193,-459,634,708,-1497,-869,2847,903,-4679,-1099,6958,2446,-9367,-7475,8549,19716,17184,8663,2663,467,36};
localparam bit [15:0] pDB19_Lo_R [38] = '{36,467,2663,8663,17184,19716,8549,-7475,-9367,2446,6958,-1099,-4679,903,2847,-869,-1497,708,634,-459,-193,230,25,-89,11,24,-9,-5,2,0,-1,0,0,-1,0,0,-1,0};
localparam bit [15:0] pDB19_Hi_D [38] = '{-37,467,-2664,8663,-17185,19716,-8550,-7475,9366,2446,-6959,-1099,4678,903,-2848,-869,1496,708,-635,-459,192,230,-26,-89,-12,24,8,-5,-3,0,0,0,-1,-1,-1,0,0,0};
localparam bit [15:0] pDB19_Hi_R [38] = '{0,0,0,-1,-1,-1,0,0,0,-3,-5,8,24,-12,-89,-26,230,192,-459,-635,708,1496,-869,-2848,903,4678,-1099,-6959,2446,9366,-7475,-8550,19716,-17185,8663,-2664,467,-37};

localparam bit [15:0] pDB20_Lo_D [40] = '{-1,0,-1,0,0,-1,-1,0,-1,-2,2,3,-13,-2,45,-28,-118,144,220,-453,-289,1058,192,-2023,184,3351,-810,-5095,1305,7480,-549,-10709,-4562,11845,20004,15489,7207,2078,345,25};
localparam bit [15:0] pDB20_Lo_R [40] = '{25,345,2078,7207,15489,20004,11845,-4562,-10709,-549,7480,1305,-5095,-810,3351,184,-2023,192,1058,-289,-453,220,144,-118,-28,45,-2,-13,3,2,-2,-1,0,-1,-1,0,0,-1,0,-1};
localparam bit [15:0] pDB20_Hi_D [40] = '{-26,345,-2079,7207,-15490,20004,-11846,-4562,10708,-549,-7481,1305,5094,-810,-3352,184,2022,192,-1059,-289,452,220,-145,-118,27,45,1,-13,-4,2,1,-1,-1,-1,0,0,-1,-1,-1,-1};
localparam bit [15:0] pDB20_Hi_R [40] = '{-1,-1,-1,-1,0,0,-1,-1,-1,1,2,-4,-13,1,45,27,-118,-145,220,452,-289,-1059,192,2022,184,-3352,-810,5094,1305,-7481,-549,10708,-4562,-11846,20004,-15490,7207,-2079,345,-26};

localparam bit [15:0] pCOIF1_Lo_D [6] = '{-514,-2384,12611,27937,11072,-2384};
localparam bit [15:0] pCOIF1_Lo_R [6] = '{-2384,11072,27937,12611,-2384,-514};
localparam bit [15:0] pCOIF1_Hi_D [6] = '{2383,11072,-27938,12611,2383,-514};
localparam bit [15:0] pCOIF1_Hi_R [6] = '{-514,2383,12611,-27938,11072,2383};

localparam bit [15:0] pCOIF2_Lo_D [12] = '{-24,-60,183,775,-1948,-2507,13664,26631,12652,-2208,-1359,536};
localparam bit [15:0] pCOIF2_Lo_R [12] = '{536,-1359,-2208,12652,26631,13664,-2507,-1948,775,183,-60,-24};
localparam bit [15:0] pCOIF2_Hi_D [12] = '{-537,-1359,2207,12652,-26632,13664,2506,-1948,-776,183,59,-24};
localparam bit [15:0] pCOIF2_Hi_R [12] = '{-24,59,183,-776,-1948,2506,13664,-26632,12652,2207,-1359,-537};

localparam bit [15:0] pCOIF3_Lo_D [18] = '{-2,-3,15,36,-85,-296,520,1132,-2697,-2353,14040,26010,13276,-2003,-2156,768,255,-125};
localparam bit [15:0] pCOIF3_Lo_R [18] = '{-125,255,768,-2156,-2003,13276,26010,14040,-2353,-2697,1132,520,-296,-85,36,15,-3,-2};
localparam bit [15:0] pCOIF3_Hi_D [18] = '{124,255,-769,-2156,2002,13276,-26011,14040,2352,-2697,-1133,520,295,-85,-37,15,2,-2};
localparam bit [15:0] pCOIF3_Hi_R [18] = '{-2,2,15,-37,-85,295,520,-1133,-2697,2352,14040,-26011,13276,2002,-2156,-769,255,124};

localparam bit [15:0] pCOIF4_Lo_D [24] = '{-1,-1,1,2,-9,-20,41,122,-186,-499,821,1288,-3153,-2184,14233,25632,13608,-1838,-2663,874,526,-241,-54,29};
localparam bit [15:0] pCOIF4_Lo_R [24] = '{29,-54,-241,526,874,-2663,-1838,13608,25632,14233,-2184,-3153,1288,821,-499,-186,122,41,-20,-9,2,1,-1,-1};
localparam bit [15:0] pCOIF4_Hi_D [24] = '{-30,-54,240,526,-875,-2663,1837,13608,-25633,14233,2183,-3153,-1289,821,498,-186,-123,41,19,-9,-3,1,0,-1};
localparam bit [15:0] pCOIF4_Hi_R [24] = '{-1,0,1,-3,-9,19,41,-123,-186,498,821,-1289,-3153,2183,14233,-25633,13608,1837,-2663,-875,526,240,-54,-30};

localparam bit [15:0] pCOIF5_Lo_D [30] = '{-1,-1,0,0,-1,-2,4,9,-21,-55,79,221,-301,-648,1070,1352,-3460,-2033,14352,25371,13813,-1706,-3013,923,767,-332,-137,71,11,-7};
localparam bit [15:0] pCOIF5_Lo_R [30] = '{-7,11,71,-137,-332,767,923,-3013,-1706,13813,25371,14352,-2033,-3460,1352,1070,-648,-301,221,79,-55,-21,9,4,-2,-1,0,0,-1,-1};
localparam bit [15:0] pCOIF5_Hi_D [30] = '{6,11,-72,-137,331,767,-924,-3013,1705,13813,-25372,14352,2032,-3460,-1353,1070,647,-301,-222,79,54,-21,-10,4,1,-1,-1,0,0,-1};
localparam bit [15:0] pCOIF5_Hi_R [30] = '{-1,0,0,-1,-1,1,4,-10,-21,54,79,-222,-301,647,1070,-1353,-3460,2032,14352,-25372,13813,1705,-3013,-924,767,331,-137,-72,11,6};

localparam bit [15:0] pSYM2_Lo_D [4] = '{-4241,7344,27410,15825};
localparam bit [15:0] pSYM2_Lo_R [4] = '{15825,27410,7344,-4241};
localparam bit [15:0] pSYM2_Hi_D [4] = '{-15826,27410,-7345,-4241};
localparam bit [15:0] pSYM2_Hi_R [4] = '{-4241,-7345,27410,-15826};

localparam bit [15:0] pSYM3_Lo_D [6] = '{1154,-2800,-4425,15069,26440,10900};
localparam bit [15:0] pSYM3_Lo_R [6] = '{10900,26440,15069,-4425,-2800,1154};
localparam bit [15:0] pSYM3_Hi_D [6] = '{-10901,26440,-15070,-4425,2799,1154};
localparam bit [15:0] pSYM3_Hi_R [6] = '{1154,2799,-4425,-15070,26440,-10901};

localparam bit [15:0] pSYM4_Lo_D [8] = '{-2483,-972,16305,26336,9760,-3252,-414,1055};
localparam bit [15:0] pSYM4_Lo_R [8] = '{1055,-414,-3252,9760,26336,16305,-972,-2483};
localparam bit [15:0] pSYM4_Hi_D [8] = '{-1056,-414,3251,9760,-26337,16305,971,-2483};
localparam bit [15:0] pSYM4_Hi_R [8] = '{-2483,971,16305,-26337,9760,3251,-414,-1056};

localparam bit [15:0] pSYM5_Lo_D [10] = '{895,967,-1283,6533,23704,20774,544,-5746,-692,640};
localparam bit [15:0] pSYM5_Lo_R [10] = '{640,-692,-5746,544,20774,23704,6533,-1283,967,895};
localparam bit [15:0] pSYM5_Hi_D [10] = '{-641,-692,5745,544,-20775,23704,-6534,-1283,-968,895};
localparam bit [15:0] pSYM5_Hi_R [10] = '{895,-968,-1283,-6534,23704,-20775,544,5745,-692,-641};

localparam bit [15:0] pSYM6_Lo_D [12] = '{504,114,-3867,-1584,16090,25809,11073,-2381,-691,1465,57,-256};
localparam bit [15:0] pSYM6_Lo_R [12] = '{-256,57,1465,-691,-2381,11073,25809,16090,-1584,-3867,114,504};
localparam bit [15:0] pSYM6_Hi_D [12] = '{255,57,-1466,-691,2380,11073,-25810,16090,1583,-3867,-115,504};
localparam bit [15:0] pSYM6_Hi_R [12] = '{504,-115,-3867,1583,16090,-25810,11073,2380,-691,-1466,57,255};

localparam bit [15:0] pSYM7_Lo_D [14] = '{87,-35,-415,999,2224,-1624,571,17566,25158,9457,-4590,-3533,131,336};
localparam bit [15:0] pSYM7_Lo_R [14] = '{336,131,-3533,-4590,9457,25158,17566,571,-1624,2224,999,-415,-35,87};
localparam bit [15:0] pSYM7_Hi_D [14] = '{-337,131,3532,-4590,-9458,25158,-17567,571,1623,2224,-1000,-415,34,87};
localparam bit [15:0] pSYM7_Hi_R [14] = '{87,34,-415,-1000,2224,1623,571,-17567,25158,-9458,-4590,3532,131,-337};

localparam bit [15:0] pSYM8_Lo_D [16] = '{-111,-18,1038,249,-4696,-2008,15773,25466,11942,-1703,-892,1610,124,-490,-10,61};
localparam bit [15:0] pSYM8_Lo_R [16] = '{61,-10,-490,124,1610,-892,-1703,11942,25466,15773,-2008,-4696,249,1038,-18,-111};
localparam bit [15:0] pSYM8_Hi_D [16] = '{-62,-10,489,124,-1611,-892,1702,11942,-25467,15773,2007,-4696,-250,1038,17,-111};
localparam bit [15:0] pSYM8_Hi_R [16] = '{-111,17,1038,-250,-4696,2007,15773,-25467,11942,1702,-892,-1611,124,489,-10,-62};

localparam bit [15:0] pSYM9_Lo_D [18] = '{45,20,-435,-378,990,19,-1789,7823,23524,20228,1155,-6277,-598,2034,290,-337,-16,35};
localparam bit [15:0] pSYM9_Lo_R [18] = '{35,-16,-337,290,2034,-598,-6277,1155,20228,23524,7823,-1789,19,990,-378,-435,20,45};
localparam bit [15:0] pSYM9_Hi_D [18] = '{-36,-16,336,290,-2035,-598,6276,1155,-20229,23524,-7824,-1789,-20,990,377,-435,-21,45};
localparam bit [15:0] pSYM9_Hi_R [18] = '{45,-21,-435,377,990,-20,-1789,-7824,23524,-20229,1155,6276,-598,-2035,290,336,-16,-36};

localparam bit [15:0] pSYM10_Lo_D [20] = '{25,3,-284,-49,1504,380,-5227,-2323,15456,25215,12577,-1165,-1049,1638,188,-667,-27,150,1,-16};
localparam bit [15:0] pSYM10_Lo_R [20] = '{-16,1,150,-27,-667,188,1638,-1049,-1165,12577,25215,15456,-2323,-5227,380,1504,-49,-284,3,25};
localparam bit [15:0] pSYM10_Hi_D [20] = '{15,1,-151,-27,666,188,-1639,-1049,1164,12577,-25216,15456,2322,-5227,-381,1504,48,-284,-4,25};
localparam bit [15:0] pSYM10_Hi_R [20] = '{25,-4,-284,48,1504,-381,-5227,2322,15456,-25216,12577,1164,-1049,-1639,188,666,-27,-151,1,15};

localparam bit [15:0] pSYM11_Lo_D [22] = '{5,-2,-57,19,213,-324,-790,1213,2292,-749,3184,18744,23931,7788,-6707,-4739,1155,1409,-66,-210,3,16};
localparam bit [15:0] pSYM11_Lo_R [22] = '{16,3,-210,-66,1409,1155,-4739,-6707,7788,23931,18744,3184,-749,2292,1213,-790,-324,213,19,-57,-2,5};
localparam bit [15:0] pSYM11_Hi_D [22] = '{-17,3,209,-66,-1410,1155,4738,-6707,-7789,23931,-18745,3184,748,2292,-1214,-790,323,213,-20,-57,1,5};
localparam bit [15:0] pSYM11_Hi_R [22] = '{5,1,-57,-20,213,323,-790,-1214,2292,748,3184,-18745,23931,-7789,-6707,4738,1155,-1410,-66,209,3,-17};

localparam bit [15:0] pSYM12_Lo_D [24] = '{3,-1,-45,5,242,-47,-794,247,1611,-1175,-727,13070,25017,15163,-2567,-5583,501,1894,-86,-479,10,77,-1,-6};
localparam bit [15:0] pSYM12_Lo_R [24] = '{-6,-1,77,10,-479,-86,1894,501,-5583,-2567,15163,25017,13070,-727,-1175,1611,247,-794,-47,242,5,-45,-1,3};
localparam bit [15:0] pSYM12_Hi_D [24] = '{5,-1,-78,10,478,-86,-1895,501,5582,-2567,-15164,25017,-13071,-727,1174,1611,-248,-794,46,242,-6,-45,0,3};
localparam bit [15:0] pSYM12_Hi_R [24] = '{3,0,-45,-6,242,46,-794,-248,1611,1174,-727,-13071,25017,-15164,-2567,5582,501,-1895,-86,478,10,-78,-1,5};

localparam bit [15:0] pSYM13_Lo_D [26] = '{2,-2,-38,-6,246,173,-663,-564,454,-1958,-4076,6478,22797,21121,3612,-4604,289,3045,577,-680,-49,185,13,-24,1,2};
localparam bit [15:0] pSYM13_Lo_R [26] = '{2,1,-24,13,185,-49,-680,577,3045,289,-4604,3612,21121,22797,6478,-4076,-1958,454,-564,-663,173,246,-6,-38,-2,2};
localparam bit [15:0] pSYM13_Hi_D [26] = '{-3,1,23,13,-186,-49,679,577,-3046,289,4603,3612,-21122,22797,-6479,-4076,1957,454,563,-663,-174,246,5,-38,1,2};
localparam bit [15:0] pSYM13_Hi_R [26] = '{2,1,-38,5,246,-174,-663,563,454,1957,-4076,-6479,22797,-21122,3612,4603,289,-3046,577,679,-49,-186,13,23,1,-3};

localparam bit [15:0] pSYM14_Lo_D [28] = '{-1,0,13,-3,-85,12,328,-91,-957,140,1226,-1889,-1158,12884,24902,15575,-1905,-5243,848,2288,-78,-637,33,148,-3,-20,0,1};
localparam bit [15:0] pSYM14_Lo_R [28] = '{1,0,-20,-3,148,33,-637,-78,2288,848,-5243,-1905,15575,24902,12884,-1158,-1889,1226,140,-957,-91,328,12,-85,-3,13,0,-1};
localparam bit [15:0] pSYM14_Hi_D [28] = '{-2,0,19,-3,-149,33,636,-78,-2289,848,5242,-1905,-15576,24902,-12885,-1158,1888,1226,-141,-957,90,328,-13,-85,2,13,-1,-1};
localparam bit [15:0] pSYM14_Hi_R [28] = '{-1,-1,13,2,-85,-13,328,90,-957,-141,1226,1888,-1158,-12885,24902,-15576,-1905,5242,848,-2289,-78,636,33,-149,-3,19,0,-2};

localparam bit [15:0] pSYM15_Lo_D [30] = '{0,-1,-6,1,35,-9,-118,112,330,-636,-1274,718,1334,-1347,3654,18960,23653,7994,-6444,-4393,2241,2227,-287,-563,50,114,-4,-14,0,0};
localparam bit [15:0] pSYM15_Lo_R [30] = '{0,0,-14,-4,114,50,-563,-287,2227,2241,-4393,-6444,7994,23653,18960,3654,-1347,1334,718,-1274,-636,330,112,-118,-9,35,1,-6,-1,0};
localparam bit [15:0] pSYM15_Hi_D [30] = '{-1,0,13,-4,-115,50,562,-287,-2228,2241,4392,-6444,-7995,23653,-18961,3654,1346,1334,-719,-1274,635,330,-113,-118,8,35,-2,-6,0,0};
localparam bit [15:0] pSYM15_Hi_R [30] = '{0,0,-6,-2,35,8,-118,-113,330,635,-1274,-719,1334,1346,3654,-18961,23653,-7995,-6444,4392,2241,-2228,-287,562,50,-115,-4,13,0,-1};

localparam bit [15:0] pSYM16_Lo_D [32] = '{0,-1,-4,0,27,-4,-128,23,415,-103,-1018,159,1059,-2195,-1133,13012,24789,15576,-1771,-5230,1006,2557,-116,-818,44,227,-8,-44,1,5,-1,-1};
localparam bit [15:0] pSYM16_Lo_R [32] = '{-1,-1,5,1,-44,-8,227,44,-818,-116,2557,1006,-5230,-1771,15576,24789,13012,-1133,-2195,1059,159,-1018,-103,415,23,-128,-4,27,0,-4,-1,0};
localparam bit [15:0] pSYM16_Hi_D [32] = '{0,-1,-6,1,43,-8,-228,44,817,-116,-2558,1006,5229,-1771,-15577,24789,-13013,-1133,2194,1059,-160,-1018,102,415,-24,-128,3,27,-1,-4,0,0};
localparam bit [15:0] pSYM16_Hi_R [32] = '{0,0,-4,-1,27,3,-128,-24,415,102,-1018,-160,1059,2194,-1133,-13013,24789,-15577,-1771,5229,1006,-2558,-116,817,44,-228,-8,43,1,-6,-1,0};

localparam bit [15:0] pSYM17_Lo_D [34] = '{0,0,-3,-1,15,-5,-90,28,343,-158,-1091,586,3432,565,-3886,4666,21322,22331,5915,-5082,-2821,529,-238,-592,326,406,-63,-129,1,23,0,-3,-1,0};
localparam bit [15:0] pSYM17_Lo_R [34] = '{0,-1,-3,0,23,1,-129,-63,406,326,-592,-238,529,-2821,-5082,5915,22331,21322,4666,-3886,565,3432,586,-1091,-158,343,28,-90,-5,15,-1,-3,0,0};
localparam bit [15:0] pSYM17_Hi_D [34] = '{-1,-1,2,0,-24,1,128,-63,-407,326,591,-238,-530,-2821,5081,5915,-22332,21322,-4667,-3886,-566,3432,-587,-1091,157,343,-29,-90,4,15,0,-3,-1,0};
localparam bit [15:0] pSYM17_Hi_R [34] = '{0,-1,-3,0,15,4,-90,-29,343,157,-1091,-587,3432,-566,-3886,-4667,21322,-22332,5915,5081,-2821,-530,-238,591,326,-407,-63,128,1,-24,0,2,-1,-1};

localparam bit [15:0] pSYM18_Lo_D [36] = '{0,0,-2,-1,12,2,-76,-14,311,53,-994,-167,2759,1113,-5241,-1705,15531,24694,13155,-1065,-2419,934,205,-1040,-107,491,35,-172,-7,46,1,-9,-1,0,0,-1};
localparam bit [15:0] pSYM18_Lo_R [36] = '{-1,0,0,-1,-9,1,46,-7,-172,35,491,-107,-1040,205,934,-2419,-1065,13155,24694,15531,-1705,-5241,1113,2759,-167,-994,53,311,-14,-76,2,12,-1,-2,0,0};
localparam bit [15:0] pSYM18_Hi_D [36] = '{0,0,-1,-1,8,1,-47,-7,171,35,-492,-107,1039,205,-935,-2419,1064,13155,-24695,15531,1704,-5241,-1114,2759,166,-994,-54,311,13,-76,-3,12,0,-2,-1,0};
localparam bit [15:0] pSYM18_Hi_R [36] = '{0,-1,-2,0,12,-3,-76,13,311,-54,-994,166,2759,-1114,-5241,1704,15531,-24695,13155,1064,-2419,-935,205,1039,-107,-492,35,171,-7,-47,1,8,-1,-1,0,0};

localparam bit [15:0] pSYM19_Lo_D [38] = '{0,-1,-1,0,3,-2,-21,5,69,-39,-168,261,517,-743,-1529,229,293,-2213,3572,18944,23578,8462,-5787,-3810,3068,2754,-555,-908,141,270,-21,-56,4,9,-1,-1,0,0};
localparam bit [15:0] pSYM19_Lo_R [38] = '{0,0,-1,-1,9,4,-56,-21,270,141,-908,-555,2754,3068,-3810,-5787,8462,23578,18944,3572,-2213,293,229,-1529,-743,517,261,-168,-39,69,5,-21,-2,3,0,-1,-1,0};
localparam bit [15:0] pSYM19_Hi_D [38] = '{-1,0,0,-1,-10,4,55,-21,-271,141,907,-555,-2755,3068,3809,-5787,-8463,23578,-18945,3572,2212,293,-230,-1529,742,517,-262,-168,38,69,-6,-21,1,3,-1,-1,0,0};
localparam bit [15:0] pSYM19_Hi_R [38] = '{0,0,-1,-1,3,1,-21,-6,69,38,-168,-262,517,742,-1529,-230,293,2212,3572,-18945,23578,-8463,-5787,3809,3068,-2755,-555,907,141,-271,-21,55,4,-10,-1,0,0,-1};

localparam bit [15:0] pSYM20_Lo_D [40] = '{0,-1,-1,0,2,-1,-17,2,68,-11,-217,46,557,-109,-1037,266,838,-2589,-978,13298,24614,15466,-1675,-5262,1187,2913,-225,-1160,63,398,-21,-114,4,24,-1,-4,0,0,-1,-1};
localparam bit [15:0] pSYM20_Lo_R [40] = '{-1,-1,0,0,-4,-1,24,4,-114,-21,398,63,-1160,-225,2913,1187,-5262,-1675,15466,24614,13298,-978,-2589,838,266,-1037,-109,557,46,-217,-11,68,2,-17,-1,2,0,-1,-1,0};
localparam bit [15:0] pSYM20_Hi_D [40] = '{0,-1,-1,0,3,-1,-25,4,113,-21,-399,63,1159,-225,-2914,1187,5261,-1675,-15467,24614,-13299,-978,2588,838,-267,-1037,108,557,-47,-217,10,68,-3,-17,0,2,-1,-1,0,0};
localparam bit [15:0] pSYM20_Hi_R [40] = '{0,0,-1,-1,2,0,-17,-3,68,10,-217,-47,557,108,-1037,-267,838,2588,-978,-13299,24614,-15467,-1675,5261,1187,-2914,-225,1159,63,-399,-21,113,4,-25,-1,3,0,-1,-1,0};

localparam bit [15:0] pDMEY_Lo_D [102] = '{0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-2,1,1,-4,0,4,-3,-5,-4,5,28,-19,-89,71,198,-210,-362,499,570,-1052,-797,2086,1003,-4349,-1149,14552,24371,14552,-1149,-4349,1003,2086,-797,-1052,570,499,-362,-210,198,71,-89,-19,28,5,-4,-5,-3,4,0,-4,1,1,-2,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1};
localparam bit [15:0] pDMEY_Lo_R [102] = '{-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-2,1,1,-4,0,4,-3,-5,-4,5,28,-19,-89,71,198,-210,-362,499,570,-1052,-797,2086,1003,-4349,-1149,14552,24371,14552,-1149,-4349,1003,2086,-797,-1052,570,499,-362,-210,198,71,-89,-19,28,5,-4,-5,-3,4,0,-4,1,1,-2,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0};
localparam bit [15:0] pDMEY_Hi_D [102] = '{0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,1,1,-2,-4,-1,4,2,-5,3,5,-29,-19,88,71,-199,-210,361,499,-571,-1052,796,2086,-1004,-4349,1148,14552,-24372,14552,1148,-4349,-1004,2086,796,-1052,-571,499,361,-210,-199,71,88,-19,-29,5,3,-5,2,4,-1,-4,-2,1,1,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0};
localparam bit [15:0] pDMEY_Hi_R [102] = '{0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,1,1,-2,-4,-1,4,2,-5,3,5,-29,-19,88,71,-199,-210,361,499,-571,-1052,796,2086,-1004,-4349,1148,14552,-24372,14552,1148,-4349,-1004,2086,796,-1052,-571,499,361,-210,-199,71,88,-19,-29,5,3,-5,2,4,-1,-4,-2,1,1,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0,0,-1,-1,-1,0,0};

